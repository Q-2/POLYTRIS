module scoreToDecimal(
    input logic [9:0]score,
    output logic [3:0]first_addr, second_addr, third_addr, fourth_addr
);
always_comb begin
unique case(score)

 10'b0: begin
first_addr = 4'h0; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101: begin
first_addr = 4'h5; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110: begin
first_addr = 4'h6; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111: begin
first_addr = 4'h7; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1000: begin
first_addr = 4'h8; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1001: begin
first_addr = 4'h9; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1010: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1011: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1100: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1101: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1110: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1111: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10000: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10001: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10010: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10011: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10100: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10101: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10110: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10111: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11000: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11001: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11010: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11011: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11100: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11101: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11110: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11111: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100000: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100001: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100010: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100011: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100100: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100101: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100110: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100111: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101000: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101001: begin
first_addr = 4'h4; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101010: begin
first_addr = 4'h4; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101011: begin
first_addr = 4'h4; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101100: begin
first_addr = 4'h4; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101101: begin
first_addr = 4'h4; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101110: begin
first_addr = 4'h4; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101111: begin
first_addr = 4'h4; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110000: begin
first_addr = 4'h4; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110001: begin
first_addr = 4'h4; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110010: begin
first_addr = 4'h5; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110011: begin
first_addr = 4'h5; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110100: begin
first_addr = 4'h5; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110101: begin
first_addr = 4'h5; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110110: begin
first_addr = 4'h5; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110111: begin
first_addr = 4'h5; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111000: begin
first_addr = 4'h5; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111001: begin
first_addr = 4'h5; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111010: begin
first_addr = 4'h5; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111011: begin
first_addr = 4'h5; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111100: begin
first_addr = 4'h6; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111101: begin
first_addr = 4'h6; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111110: begin
first_addr = 4'h6; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111111: begin
first_addr = 4'h6; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1000000: begin
first_addr = 4'h6; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1000001: begin
first_addr = 4'h6; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1000010: begin
first_addr = 4'h6; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1000011: begin
first_addr = 4'h6; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1000100: begin
first_addr = 4'h6; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1000101: begin
first_addr = 4'h6; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1000110: begin
first_addr = 4'h7; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1000111: begin
first_addr = 4'h7; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1001000: begin
first_addr = 4'h7; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1001001: begin
first_addr = 4'h7; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1001010: begin
first_addr = 4'h7; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1001011: begin
first_addr = 4'h7; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1001100: begin
first_addr = 4'h7; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1001101: begin
first_addr = 4'h7; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1001110: begin
first_addr = 4'h7; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1001111: begin
first_addr = 4'h7; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1010000: begin
first_addr = 4'h8; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1010001: begin
first_addr = 4'h8; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1010010: begin
first_addr = 4'h8; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1010011: begin
first_addr = 4'h8; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1010100: begin
first_addr = 4'h8; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1010101: begin
first_addr = 4'h8; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1010110: begin
first_addr = 4'h8; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1010111: begin
first_addr = 4'h8; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1011000: begin
first_addr = 4'h8; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1011001: begin
first_addr = 4'h8; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1011010: begin
first_addr = 4'h9; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1011011: begin
first_addr = 4'h9; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1011100: begin
first_addr = 4'h9; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1011101: begin
first_addr = 4'h9; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1011110: begin
first_addr = 4'h9; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1011111: begin
first_addr = 4'h9; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1100000: begin
first_addr = 4'h9; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1100001: begin
first_addr = 4'h9; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1100010: begin
first_addr = 4'h9; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1100011: begin
first_addr = 4'h9; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1100100: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1100101: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1100110: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1100111: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1101000: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1101001: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1101010: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1101011: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1101100: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1101101: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1101110: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1101111: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1110000: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1110001: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1110010: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1110011: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1110100: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1110101: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1110110: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1110111: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1111000: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1111001: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1111010: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1111011: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1111100: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1111101: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1111110: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1111111: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b10000000: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b10000001: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b10000010: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10000011: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b10000100: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b10000101: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b10000110: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b10000111: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b10001000: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b10001001: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b10001010: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b10001011: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b10001100: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10001101: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b10001110: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b10001111: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b10010000: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b10010001: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b10010010: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b10010011: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b10010100: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b10010101: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b10010110: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10010111: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b10011000: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b10011001: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b10011010: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b10011011: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b10011100: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b10011101: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b10011110: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b10011111: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b10100000: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10100001: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b10100010: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b10100011: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b10100100: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b10100101: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b10100110: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b10100111: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b10101000: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b10101001: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b10101010: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10101011: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b10101100: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b10101101: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b10101110: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b10101111: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b10110000: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b10110001: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b10110010: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b10110011: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b10110100: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10110101: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b10110110: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b10110111: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b10111000: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b10111001: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b10111010: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b10111011: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b10111100: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b10111101: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b10111110: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10111111: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b11000000: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b11000001: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b11000010: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b11000011: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b11000100: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b11000101: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b11000110: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b11000111: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b11001000: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11001001: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b11001010: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b11001011: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b11001100: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b11001101: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b11001110: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b11001111: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b11010000: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b11010001: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b11010010: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11010011: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b11010100: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b11010101: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b11010110: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b11010111: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b11011000: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b11011001: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b11011010: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b11011011: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b11011100: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11011101: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b11011110: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b11011111: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b11100000: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b11100001: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b11100010: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b11100011: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b11100100: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b11100101: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b11100110: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11100111: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b11101000: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b11101001: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b11101010: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b11101011: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b11101100: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b11101101: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b11101110: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b11101111: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b11110000: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11110001: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b11110010: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b11110011: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b11110100: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b11110101: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b11110110: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b11110111: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b11111000: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b11111001: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b11111010: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11111011: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b11111100: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b11111101: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b11111110: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b11111111: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b100000000: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b100000001: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b100000010: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b100000011: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b100000100: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100000101: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b100000110: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b100000111: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b100001000: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b100001001: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b100001010: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b100001011: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b100001100: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b100001101: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b100001110: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100001111: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b100010000: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b100010001: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b100010010: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b100010011: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b100010100: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b100010101: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b100010110: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b100010111: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b100011000: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100011001: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b100011010: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b100011011: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b100011100: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b100011101: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b100011110: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b100011111: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b100100000: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b100100001: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b100100010: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100100011: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b100100100: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b100100101: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b100100110: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b100100111: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b100101000: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b100101001: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b100101010: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b100101011: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b100101100: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100101101: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b100101110: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b100101111: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b100110000: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b100110001: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b100110010: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b100110011: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b100110100: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b100110101: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b100110110: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100110111: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b100111000: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b100111001: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b100111010: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b100111011: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b100111100: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b100111101: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b100111110: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b100111111: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b101000000: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101000001: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b101000010: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b101000011: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b101000100: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b101000101: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b101000110: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b101000111: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b101001000: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b101001001: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b101001010: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101001011: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b101001100: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b101001101: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b101001110: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b101001111: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b101010000: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b101010001: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b101010010: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b101010011: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b101010100: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101010101: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b101010110: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b101010111: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b101011000: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b101011001: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b101011010: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b101011011: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b101011100: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b101011101: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b101011110: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101011111: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b101100000: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b101100001: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b101100010: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b101100011: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b101100100: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b101100101: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b101100110: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b101100111: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b101101000: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101101001: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b101101010: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b101101011: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b101101100: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b101101101: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b101101110: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b101101111: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b101110000: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b101110001: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b101110010: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101110011: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b101110100: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b101110101: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b101110110: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b101110111: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b101111000: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b101111001: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b101111010: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b101111011: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b101111100: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101111101: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b101111110: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b101111111: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b110000000: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b110000001: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b110000010: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b110000011: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b110000100: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b110000101: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b110000110: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110000111: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b110001000: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b110001001: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b110001010: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b110001011: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b110001100: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b110001101: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b110001110: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b110001111: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b110010000: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110010001: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b110010010: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b110010011: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b110010100: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b110010101: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b110010110: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b110010111: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b110011000: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b110011001: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b110011010: begin
first_addr = 4'h4; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110011011: begin
first_addr = 4'h4; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b110011100: begin
first_addr = 4'h4; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b110011101: begin
first_addr = 4'h4; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b110011110: begin
first_addr = 4'h4; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b110011111: begin
first_addr = 4'h4; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b110100000: begin
first_addr = 4'h4; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b110100001: begin
first_addr = 4'h4; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b110100010: begin
first_addr = 4'h4; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b110100011: begin
first_addr = 4'h4; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b110100100: begin
first_addr = 4'h4; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110100101: begin
first_addr = 4'h4; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b110100110: begin
first_addr = 4'h4; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b110100111: begin
first_addr = 4'h4; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b110101000: begin
first_addr = 4'h4; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b110101001: begin
first_addr = 4'h4; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b110101010: begin
first_addr = 4'h4; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b110101011: begin
first_addr = 4'h4; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b110101100: begin
first_addr = 4'h4; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b110101101: begin
first_addr = 4'h4; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b110101110: begin
first_addr = 4'h4; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110101111: begin
first_addr = 4'h4; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b110110000: begin
first_addr = 4'h4; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b110110001: begin
first_addr = 4'h4; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b110110010: begin
first_addr = 4'h4; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b110110011: begin
first_addr = 4'h4; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b110110100: begin
first_addr = 4'h4; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b110110101: begin
first_addr = 4'h4; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b110110110: begin
first_addr = 4'h4; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b110110111: begin
first_addr = 4'h4; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b110111000: begin
first_addr = 4'h4; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110111001: begin
first_addr = 4'h4; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b110111010: begin
first_addr = 4'h4; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b110111011: begin
first_addr = 4'h4; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b110111100: begin
first_addr = 4'h4; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b110111101: begin
first_addr = 4'h4; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b110111110: begin
first_addr = 4'h4; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b110111111: begin
first_addr = 4'h4; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b111000000: begin
first_addr = 4'h4; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b111000001: begin
first_addr = 4'h4; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b111000010: begin
first_addr = 4'h4; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111000011: begin
first_addr = 4'h4; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b111000100: begin
first_addr = 4'h4; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b111000101: begin
first_addr = 4'h4; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b111000110: begin
first_addr = 4'h4; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b111000111: begin
first_addr = 4'h4; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b111001000: begin
first_addr = 4'h4; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b111001001: begin
first_addr = 4'h4; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b111001010: begin
first_addr = 4'h4; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b111001011: begin
first_addr = 4'h4; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b111001100: begin
first_addr = 4'h4; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111001101: begin
first_addr = 4'h4; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b111001110: begin
first_addr = 4'h4; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b111001111: begin
first_addr = 4'h4; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b111010000: begin
first_addr = 4'h4; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b111010001: begin
first_addr = 4'h4; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b111010010: begin
first_addr = 4'h4; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b111010011: begin
first_addr = 4'h4; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b111010100: begin
first_addr = 4'h4; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b111010101: begin
first_addr = 4'h4; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b111010110: begin
first_addr = 4'h4; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111010111: begin
first_addr = 4'h4; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b111011000: begin
first_addr = 4'h4; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b111011001: begin
first_addr = 4'h4; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b111011010: begin
first_addr = 4'h4; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b111011011: begin
first_addr = 4'h4; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b111011100: begin
first_addr = 4'h4; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b111011101: begin
first_addr = 4'h4; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b111011110: begin
first_addr = 4'h4; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b111011111: begin
first_addr = 4'h4; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b111100000: begin
first_addr = 4'h4; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111100001: begin
first_addr = 4'h4; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b111100010: begin
first_addr = 4'h4; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b111100011: begin
first_addr = 4'h4; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b111100100: begin
first_addr = 4'h4; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b111100101: begin
first_addr = 4'h4; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b111100110: begin
first_addr = 4'h4; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b111100111: begin
first_addr = 4'h4; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b111101000: begin
first_addr = 4'h4; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b111101001: begin
first_addr = 4'h4; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b111101010: begin
first_addr = 4'h4; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111101011: begin
first_addr = 4'h4; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b111101100: begin
first_addr = 4'h4; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b111101101: begin
first_addr = 4'h4; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b111101110: begin
first_addr = 4'h4; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b111101111: begin
first_addr = 4'h4; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b111110000: begin
first_addr = 4'h4; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b111110001: begin
first_addr = 4'h4; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b111110010: begin
first_addr = 4'h4; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b111110011: begin
first_addr = 4'h4; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b111110100: begin
first_addr = 4'h5; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111110101: begin
first_addr = 4'h5; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b111110110: begin
first_addr = 4'h5; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b111110111: begin
first_addr = 4'h5; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b111111000: begin
first_addr = 4'h5; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b111111001: begin
first_addr = 4'h5; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b111111010: begin
first_addr = 4'h5; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b111111011: begin
first_addr = 4'h5; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b111111100: begin
first_addr = 4'h5; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b111111101: begin
first_addr = 4'h5; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b111111110: begin
first_addr = 4'h5; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111111111: begin
first_addr = 4'h5; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1000000000: begin
first_addr = 4'h5; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1000000001: begin
first_addr = 4'h5; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1000000010: begin
first_addr = 4'h5; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1000000011: begin
first_addr = 4'h5; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1000000100: begin
first_addr = 4'h5; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1000000101: begin
first_addr = 4'h5; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1000000110: begin
first_addr = 4'h5; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1000000111: begin
first_addr = 4'h5; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1000001000: begin
first_addr = 4'h5; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1000001001: begin
first_addr = 4'h5; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1000001010: begin
first_addr = 4'h5; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1000001011: begin
first_addr = 4'h5; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1000001100: begin
first_addr = 4'h5; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1000001101: begin
first_addr = 4'h5; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1000001110: begin
first_addr = 4'h5; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1000001111: begin
first_addr = 4'h5; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1000010000: begin
first_addr = 4'h5; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1000010001: begin
first_addr = 4'h5; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1000010010: begin
first_addr = 4'h5; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1000010011: begin
first_addr = 4'h5; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1000010100: begin
first_addr = 4'h5; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1000010101: begin
first_addr = 4'h5; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1000010110: begin
first_addr = 4'h5; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1000010111: begin
first_addr = 4'h5; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1000011000: begin
first_addr = 4'h5; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1000011001: begin
first_addr = 4'h5; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1000011010: begin
first_addr = 4'h5; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1000011011: begin
first_addr = 4'h5; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1000011100: begin
first_addr = 4'h5; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1000011101: begin
first_addr = 4'h5; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1000011110: begin
first_addr = 4'h5; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1000011111: begin
first_addr = 4'h5; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1000100000: begin
first_addr = 4'h5; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1000100001: begin
first_addr = 4'h5; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1000100010: begin
first_addr = 4'h5; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1000100011: begin
first_addr = 4'h5; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1000100100: begin
first_addr = 4'h5; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1000100101: begin
first_addr = 4'h5; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1000100110: begin
first_addr = 4'h5; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1000100111: begin
first_addr = 4'h5; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1000101000: begin
first_addr = 4'h5; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1000101001: begin
first_addr = 4'h5; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1000101010: begin
first_addr = 4'h5; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1000101011: begin
first_addr = 4'h5; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1000101100: begin
first_addr = 4'h5; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1000101101: begin
first_addr = 4'h5; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1000101110: begin
first_addr = 4'h5; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1000101111: begin
first_addr = 4'h5; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1000110000: begin
first_addr = 4'h5; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1000110001: begin
first_addr = 4'h5; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1000110010: begin
first_addr = 4'h5; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1000110011: begin
first_addr = 4'h5; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1000110100: begin
first_addr = 4'h5; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1000110101: begin
first_addr = 4'h5; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1000110110: begin
first_addr = 4'h5; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1000110111: begin
first_addr = 4'h5; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1000111000: begin
first_addr = 4'h5; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1000111001: begin
first_addr = 4'h5; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1000111010: begin
first_addr = 4'h5; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1000111011: begin
first_addr = 4'h5; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1000111100: begin
first_addr = 4'h5; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1000111101: begin
first_addr = 4'h5; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1000111110: begin
first_addr = 4'h5; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1000111111: begin
first_addr = 4'h5; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1001000000: begin
first_addr = 4'h5; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1001000001: begin
first_addr = 4'h5; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1001000010: begin
first_addr = 4'h5; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1001000011: begin
first_addr = 4'h5; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1001000100: begin
first_addr = 4'h5; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1001000101: begin
first_addr = 4'h5; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1001000110: begin
first_addr = 4'h5; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1001000111: begin
first_addr = 4'h5; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1001001000: begin
first_addr = 4'h5; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1001001001: begin
first_addr = 4'h5; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1001001010: begin
first_addr = 4'h5; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1001001011: begin
first_addr = 4'h5; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1001001100: begin
first_addr = 4'h5; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1001001101: begin
first_addr = 4'h5; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1001001110: begin
first_addr = 4'h5; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1001001111: begin
first_addr = 4'h5; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1001010000: begin
first_addr = 4'h5; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1001010001: begin
first_addr = 4'h5; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1001010010: begin
first_addr = 4'h5; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1001010011: begin
first_addr = 4'h5; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1001010100: begin
first_addr = 4'h5; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1001010101: begin
first_addr = 4'h5; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1001010110: begin
first_addr = 4'h5; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1001010111: begin
first_addr = 4'h5; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1001011000: begin
first_addr = 4'h6; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1001011001: begin
first_addr = 4'h6; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1001011010: begin
first_addr = 4'h6; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1001011011: begin
first_addr = 4'h6; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1001011100: begin
first_addr = 4'h6; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1001011101: begin
first_addr = 4'h6; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1001011110: begin
first_addr = 4'h6; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1001011111: begin
first_addr = 4'h6; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1001100000: begin
first_addr = 4'h6; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1001100001: begin
first_addr = 4'h6; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1001100010: begin
first_addr = 4'h6; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1001100011: begin
first_addr = 4'h6; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1001100100: begin
first_addr = 4'h6; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1001100101: begin
first_addr = 4'h6; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1001100110: begin
first_addr = 4'h6; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1001100111: begin
first_addr = 4'h6; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1001101000: begin
first_addr = 4'h6; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1001101001: begin
first_addr = 4'h6; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1001101010: begin
first_addr = 4'h6; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1001101011: begin
first_addr = 4'h6; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1001101100: begin
first_addr = 4'h6; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1001101101: begin
first_addr = 4'h6; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1001101110: begin
first_addr = 4'h6; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1001101111: begin
first_addr = 4'h6; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1001110000: begin
first_addr = 4'h6; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1001110001: begin
first_addr = 4'h6; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1001110010: begin
first_addr = 4'h6; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1001110011: begin
first_addr = 4'h6; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1001110100: begin
first_addr = 4'h6; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1001110101: begin
first_addr = 4'h6; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1001110110: begin
first_addr = 4'h6; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1001110111: begin
first_addr = 4'h6; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1001111000: begin
first_addr = 4'h6; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1001111001: begin
first_addr = 4'h6; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1001111010: begin
first_addr = 4'h6; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1001111011: begin
first_addr = 4'h6; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1001111100: begin
first_addr = 4'h6; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1001111101: begin
first_addr = 4'h6; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1001111110: begin
first_addr = 4'h6; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1001111111: begin
first_addr = 4'h6; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1010000000: begin
first_addr = 4'h6; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1010000001: begin
first_addr = 4'h6; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1010000010: begin
first_addr = 4'h6; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1010000011: begin
first_addr = 4'h6; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1010000100: begin
first_addr = 4'h6; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1010000101: begin
first_addr = 4'h6; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1010000110: begin
first_addr = 4'h6; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1010000111: begin
first_addr = 4'h6; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1010001000: begin
first_addr = 4'h6; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1010001001: begin
first_addr = 4'h6; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1010001010: begin
first_addr = 4'h6; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1010001011: begin
first_addr = 4'h6; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1010001100: begin
first_addr = 4'h6; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1010001101: begin
first_addr = 4'h6; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1010001110: begin
first_addr = 4'h6; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1010001111: begin
first_addr = 4'h6; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1010010000: begin
first_addr = 4'h6; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1010010001: begin
first_addr = 4'h6; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1010010010: begin
first_addr = 4'h6; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1010010011: begin
first_addr = 4'h6; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1010010100: begin
first_addr = 4'h6; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1010010101: begin
first_addr = 4'h6; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1010010110: begin
first_addr = 4'h6; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1010010111: begin
first_addr = 4'h6; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1010011000: begin
first_addr = 4'h6; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1010011001: begin
first_addr = 4'h6; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1010011010: begin
first_addr = 4'h6; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1010011011: begin
first_addr = 4'h6; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1010011100: begin
first_addr = 4'h6; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1010011101: begin
first_addr = 4'h6; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1010011110: begin
first_addr = 4'h6; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1010011111: begin
first_addr = 4'h6; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1010100000: begin
first_addr = 4'h6; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1010100001: begin
first_addr = 4'h6; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1010100010: begin
first_addr = 4'h6; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1010100011: begin
first_addr = 4'h6; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1010100100: begin
first_addr = 4'h6; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1010100101: begin
first_addr = 4'h6; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1010100110: begin
first_addr = 4'h6; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1010100111: begin
first_addr = 4'h6; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1010101000: begin
first_addr = 4'h6; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1010101001: begin
first_addr = 4'h6; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1010101010: begin
first_addr = 4'h6; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1010101011: begin
first_addr = 4'h6; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1010101100: begin
first_addr = 4'h6; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1010101101: begin
first_addr = 4'h6; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1010101110: begin
first_addr = 4'h6; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1010101111: begin
first_addr = 4'h6; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1010110000: begin
first_addr = 4'h6; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1010110001: begin
first_addr = 4'h6; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1010110010: begin
first_addr = 4'h6; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1010110011: begin
first_addr = 4'h6; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1010110100: begin
first_addr = 4'h6; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1010110101: begin
first_addr = 4'h6; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1010110110: begin
first_addr = 4'h6; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1010110111: begin
first_addr = 4'h6; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1010111000: begin
first_addr = 4'h6; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1010111001: begin
first_addr = 4'h6; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1010111010: begin
first_addr = 4'h6; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1010111011: begin
first_addr = 4'h6; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1010111100: begin
first_addr = 4'h7; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1010111101: begin
first_addr = 4'h7; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1010111110: begin
first_addr = 4'h7; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1010111111: begin
first_addr = 4'h7; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1011000000: begin
first_addr = 4'h7; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1011000001: begin
first_addr = 4'h7; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1011000010: begin
first_addr = 4'h7; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1011000011: begin
first_addr = 4'h7; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1011000100: begin
first_addr = 4'h7; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1011000101: begin
first_addr = 4'h7; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1011000110: begin
first_addr = 4'h7; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1011000111: begin
first_addr = 4'h7; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1011001000: begin
first_addr = 4'h7; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1011001001: begin
first_addr = 4'h7; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1011001010: begin
first_addr = 4'h7; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1011001011: begin
first_addr = 4'h7; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1011001100: begin
first_addr = 4'h7; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1011001101: begin
first_addr = 4'h7; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1011001110: begin
first_addr = 4'h7; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1011001111: begin
first_addr = 4'h7; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1011010000: begin
first_addr = 4'h7; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1011010001: begin
first_addr = 4'h7; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1011010010: begin
first_addr = 4'h7; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1011010011: begin
first_addr = 4'h7; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1011010100: begin
first_addr = 4'h7; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1011010101: begin
first_addr = 4'h7; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1011010110: begin
first_addr = 4'h7; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1011010111: begin
first_addr = 4'h7; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1011011000: begin
first_addr = 4'h7; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1011011001: begin
first_addr = 4'h7; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1011011010: begin
first_addr = 4'h7; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1011011011: begin
first_addr = 4'h7; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1011011100: begin
first_addr = 4'h7; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1011011101: begin
first_addr = 4'h7; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1011011110: begin
first_addr = 4'h7; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1011011111: begin
first_addr = 4'h7; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1011100000: begin
first_addr = 4'h7; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1011100001: begin
first_addr = 4'h7; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1011100010: begin
first_addr = 4'h7; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1011100011: begin
first_addr = 4'h7; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1011100100: begin
first_addr = 4'h7; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1011100101: begin
first_addr = 4'h7; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1011100110: begin
first_addr = 4'h7; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1011100111: begin
first_addr = 4'h7; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1011101000: begin
first_addr = 4'h7; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1011101001: begin
first_addr = 4'h7; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1011101010: begin
first_addr = 4'h7; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1011101011: begin
first_addr = 4'h7; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1011101100: begin
first_addr = 4'h7; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1011101101: begin
first_addr = 4'h7; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1011101110: begin
first_addr = 4'h7; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1011101111: begin
first_addr = 4'h7; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1011110000: begin
first_addr = 4'h7; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1011110001: begin
first_addr = 4'h7; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1011110010: begin
first_addr = 4'h7; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1011110011: begin
first_addr = 4'h7; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1011110100: begin
first_addr = 4'h7; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1011110101: begin
first_addr = 4'h7; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1011110110: begin
first_addr = 4'h7; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1011110111: begin
first_addr = 4'h7; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1011111000: begin
first_addr = 4'h7; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1011111001: begin
first_addr = 4'h7; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1011111010: begin
first_addr = 4'h7; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1011111011: begin
first_addr = 4'h7; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1011111100: begin
first_addr = 4'h7; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1011111101: begin
first_addr = 4'h7; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1011111110: begin
first_addr = 4'h7; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1011111111: begin
first_addr = 4'h7; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1100000000: begin
first_addr = 4'h7; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1100000001: begin
first_addr = 4'h7; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1100000010: begin
first_addr = 4'h7; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1100000011: begin
first_addr = 4'h7; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1100000100: begin
first_addr = 4'h7; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1100000101: begin
first_addr = 4'h7; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1100000110: begin
first_addr = 4'h7; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1100000111: begin
first_addr = 4'h7; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1100001000: begin
first_addr = 4'h7; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1100001001: begin
first_addr = 4'h7; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1100001010: begin
first_addr = 4'h7; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1100001011: begin
first_addr = 4'h7; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1100001100: begin
first_addr = 4'h7; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1100001101: begin
first_addr = 4'h7; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1100001110: begin
first_addr = 4'h7; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1100001111: begin
first_addr = 4'h7; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1100010000: begin
first_addr = 4'h7; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1100010001: begin
first_addr = 4'h7; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1100010010: begin
first_addr = 4'h7; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1100010011: begin
first_addr = 4'h7; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1100010100: begin
first_addr = 4'h7; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1100010101: begin
first_addr = 4'h7; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1100010110: begin
first_addr = 4'h7; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1100010111: begin
first_addr = 4'h7; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1100011000: begin
first_addr = 4'h7; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1100011001: begin
first_addr = 4'h7; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1100011010: begin
first_addr = 4'h7; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1100011011: begin
first_addr = 4'h7; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1100011100: begin
first_addr = 4'h7; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1100011101: begin
first_addr = 4'h7; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1100011110: begin
first_addr = 4'h7; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1100011111: begin
first_addr = 4'h7; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1100100000: begin
first_addr = 4'h8; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1100100001: begin
first_addr = 4'h8; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1100100010: begin
first_addr = 4'h8; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1100100011: begin
first_addr = 4'h8; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1100100100: begin
first_addr = 4'h8; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1100100101: begin
first_addr = 4'h8; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1100100110: begin
first_addr = 4'h8; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1100100111: begin
first_addr = 4'h8; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1100101000: begin
first_addr = 4'h8; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1100101001: begin
first_addr = 4'h8; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1100101010: begin
first_addr = 4'h8; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1100101011: begin
first_addr = 4'h8; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1100101100: begin
first_addr = 4'h8; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1100101101: begin
first_addr = 4'h8; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1100101110: begin
first_addr = 4'h8; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1100101111: begin
first_addr = 4'h8; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1100110000: begin
first_addr = 4'h8; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1100110001: begin
first_addr = 4'h8; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1100110010: begin
first_addr = 4'h8; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1100110011: begin
first_addr = 4'h8; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1100110100: begin
first_addr = 4'h8; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1100110101: begin
first_addr = 4'h8; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1100110110: begin
first_addr = 4'h8; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1100110111: begin
first_addr = 4'h8; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1100111000: begin
first_addr = 4'h8; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1100111001: begin
first_addr = 4'h8; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1100111010: begin
first_addr = 4'h8; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1100111011: begin
first_addr = 4'h8; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1100111100: begin
first_addr = 4'h8; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1100111101: begin
first_addr = 4'h8; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1100111110: begin
first_addr = 4'h8; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1100111111: begin
first_addr = 4'h8; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1101000000: begin
first_addr = 4'h8; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1101000001: begin
first_addr = 4'h8; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1101000010: begin
first_addr = 4'h8; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1101000011: begin
first_addr = 4'h8; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1101000100: begin
first_addr = 4'h8; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1101000101: begin
first_addr = 4'h8; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1101000110: begin
first_addr = 4'h8; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1101000111: begin
first_addr = 4'h8; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1101001000: begin
first_addr = 4'h8; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1101001001: begin
first_addr = 4'h8; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1101001010: begin
first_addr = 4'h8; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1101001011: begin
first_addr = 4'h8; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1101001100: begin
first_addr = 4'h8; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1101001101: begin
first_addr = 4'h8; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1101001110: begin
first_addr = 4'h8; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1101001111: begin
first_addr = 4'h8; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1101010000: begin
first_addr = 4'h8; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1101010001: begin
first_addr = 4'h8; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1101010010: begin
first_addr = 4'h8; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1101010011: begin
first_addr = 4'h8; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1101010100: begin
first_addr = 4'h8; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1101010101: begin
first_addr = 4'h8; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1101010110: begin
first_addr = 4'h8; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1101010111: begin
first_addr = 4'h8; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1101011000: begin
first_addr = 4'h8; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1101011001: begin
first_addr = 4'h8; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1101011010: begin
first_addr = 4'h8; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1101011011: begin
first_addr = 4'h8; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1101011100: begin
first_addr = 4'h8; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1101011101: begin
first_addr = 4'h8; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1101011110: begin
first_addr = 4'h8; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1101011111: begin
first_addr = 4'h8; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1101100000: begin
first_addr = 4'h8; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1101100001: begin
first_addr = 4'h8; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1101100010: begin
first_addr = 4'h8; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1101100011: begin
first_addr = 4'h8; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1101100100: begin
first_addr = 4'h8; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1101100101: begin
first_addr = 4'h8; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1101100110: begin
first_addr = 4'h8; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1101100111: begin
first_addr = 4'h8; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1101101000: begin
first_addr = 4'h8; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1101101001: begin
first_addr = 4'h8; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1101101010: begin
first_addr = 4'h8; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1101101011: begin
first_addr = 4'h8; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1101101100: begin
first_addr = 4'h8; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1101101101: begin
first_addr = 4'h8; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1101101110: begin
first_addr = 4'h8; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1101101111: begin
first_addr = 4'h8; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1101110000: begin
first_addr = 4'h8; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1101110001: begin
first_addr = 4'h8; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1101110010: begin
first_addr = 4'h8; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1101110011: begin
first_addr = 4'h8; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1101110100: begin
first_addr = 4'h8; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1101110101: begin
first_addr = 4'h8; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1101110110: begin
first_addr = 4'h8; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1101110111: begin
first_addr = 4'h8; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1101111000: begin
first_addr = 4'h8; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1101111001: begin
first_addr = 4'h8; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1101111010: begin
first_addr = 4'h8; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1101111011: begin
first_addr = 4'h8; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1101111100: begin
first_addr = 4'h8; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1101111101: begin
first_addr = 4'h8; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1101111110: begin
first_addr = 4'h8; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1101111111: begin
first_addr = 4'h8; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1110000000: begin
first_addr = 4'h8; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1110000001: begin
first_addr = 4'h8; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1110000010: begin
first_addr = 4'h8; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1110000011: begin
first_addr = 4'h8; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1110000100: begin
first_addr = 4'h9; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1110000101: begin
first_addr = 4'h9; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1110000110: begin
first_addr = 4'h9; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1110000111: begin
first_addr = 4'h9; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1110001000: begin
first_addr = 4'h9; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1110001001: begin
first_addr = 4'h9; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1110001010: begin
first_addr = 4'h9; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1110001011: begin
first_addr = 4'h9; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1110001100: begin
first_addr = 4'h9; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1110001101: begin
first_addr = 4'h9; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1110001110: begin
first_addr = 4'h9; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1110001111: begin
first_addr = 4'h9; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1110010000: begin
first_addr = 4'h9; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1110010001: begin
first_addr = 4'h9; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1110010010: begin
first_addr = 4'h9; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1110010011: begin
first_addr = 4'h9; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1110010100: begin
first_addr = 4'h9; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1110010101: begin
first_addr = 4'h9; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1110010110: begin
first_addr = 4'h9; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1110010111: begin
first_addr = 4'h9; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1110011000: begin
first_addr = 4'h9; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1110011001: begin
first_addr = 4'h9; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1110011010: begin
first_addr = 4'h9; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1110011011: begin
first_addr = 4'h9; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1110011100: begin
first_addr = 4'h9; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1110011101: begin
first_addr = 4'h9; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1110011110: begin
first_addr = 4'h9; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1110011111: begin
first_addr = 4'h9; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1110100000: begin
first_addr = 4'h9; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1110100001: begin
first_addr = 4'h9; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1110100010: begin
first_addr = 4'h9; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1110100011: begin
first_addr = 4'h9; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1110100100: begin
first_addr = 4'h9; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1110100101: begin
first_addr = 4'h9; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1110100110: begin
first_addr = 4'h9; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1110100111: begin
first_addr = 4'h9; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1110101000: begin
first_addr = 4'h9; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1110101001: begin
first_addr = 4'h9; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1110101010: begin
first_addr = 4'h9; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1110101011: begin
first_addr = 4'h9; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1110101100: begin
first_addr = 4'h9; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1110101101: begin
first_addr = 4'h9; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1110101110: begin
first_addr = 4'h9; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1110101111: begin
first_addr = 4'h9; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1110110000: begin
first_addr = 4'h9; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1110110001: begin
first_addr = 4'h9; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1110110010: begin
first_addr = 4'h9; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1110110011: begin
first_addr = 4'h9; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1110110100: begin
first_addr = 4'h9; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1110110101: begin
first_addr = 4'h9; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1110110110: begin
first_addr = 4'h9; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1110110111: begin
first_addr = 4'h9; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1110111000: begin
first_addr = 4'h9; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1110111001: begin
first_addr = 4'h9; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1110111010: begin
first_addr = 4'h9; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1110111011: begin
first_addr = 4'h9; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1110111100: begin
first_addr = 4'h9; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1110111101: begin
first_addr = 4'h9; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1110111110: begin
first_addr = 4'h9; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1110111111: begin
first_addr = 4'h9; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1111000000: begin
first_addr = 4'h9; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1111000001: begin
first_addr = 4'h9; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1111000010: begin
first_addr = 4'h9; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1111000011: begin
first_addr = 4'h9; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1111000100: begin
first_addr = 4'h9; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1111000101: begin
first_addr = 4'h9; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1111000110: begin
first_addr = 4'h9; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1111000111: begin
first_addr = 4'h9; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1111001000: begin
first_addr = 4'h9; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1111001001: begin
first_addr = 4'h9; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1111001010: begin
first_addr = 4'h9; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1111001011: begin
first_addr = 4'h9; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1111001100: begin
first_addr = 4'h9; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1111001101: begin
first_addr = 4'h9; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1111001110: begin
first_addr = 4'h9; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1111001111: begin
first_addr = 4'h9; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1111010000: begin
first_addr = 4'h9; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1111010001: begin
first_addr = 4'h9; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1111010010: begin
first_addr = 4'h9; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1111010011: begin
first_addr = 4'h9; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1111010100: begin
first_addr = 4'h9; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1111010101: begin
first_addr = 4'h9; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1111010110: begin
first_addr = 4'h9; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1111010111: begin
first_addr = 4'h9; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1111011000: begin
first_addr = 4'h9; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1111011001: begin
first_addr = 4'h9; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1111011010: begin
first_addr = 4'h9; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1111011011: begin
first_addr = 4'h9; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1111011100: begin
first_addr = 4'h9; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1111011101: begin
first_addr = 4'h9; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1111011110: begin
first_addr = 4'h9; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1111011111: begin
first_addr = 4'h9; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1111100000: begin
first_addr = 4'h9; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1111100001: begin
first_addr = 4'h9; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b1111100010: begin
first_addr = 4'h9; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b1111100011: begin
first_addr = 4'h9; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b1111100100: begin
first_addr = 4'h9; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b1111100101: begin
first_addr = 4'h9; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b1111100110: begin
first_addr = 4'h9; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b1111100111: begin
first_addr = 4'h9; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b1111101000: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b1111101001: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b1111101010: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b1111101011: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b1111101100: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b1111101101: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b1111101110: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b1111101111: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b1111110000: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b1111110001: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b1111110010: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b1111110011: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b1111110100: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b1111110101: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b1111110110: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b1111110111: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b1111111000: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b1111111001: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b1111111010: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b1111111011: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b1111111100: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b1111111101: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b1111111110: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b1111111111: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b10000000000: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b10000000001: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b10000000010: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b10000000011: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b10000000100: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b10000000101: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b10000000110: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b10000000111: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b10000001000: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b10000001001: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b10000001010: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b10000001011: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b10000001100: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b10000001101: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b10000001110: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b10000001111: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b10000010000: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b10000010001: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b10000010010: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b10000010011: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b10000010100: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b10000010101: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b10000010110: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b10000010111: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b10000011000: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b10000011001: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b10000011010: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b10000011011: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b10000011100: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b10000011101: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b10000011110: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b10000011111: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b10000100000: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b10000100001: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b10000100010: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b10000100011: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b10000100100: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b10000100101: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b10000100110: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b10000100111: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b10000101000: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b10000101001: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b10000101010: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b10000101011: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b10000101100: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b10000101101: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b10000101110: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b10000101111: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b10000110000: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b10000110001: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b10000110010: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b10000110011: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b10000110100: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b10000110101: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b10000110110: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b10000110111: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b10000111000: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b10000111001: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b10000111010: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b10000111011: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b10000111100: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b10000111101: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b10000111110: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b10000111111: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b10001000000: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b10001000001: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b10001000010: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b10001000011: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b10001000100: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b10001000101: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b10001000110: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b10001000111: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b10001001000: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b10001001001: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b10001001010: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b10001001011: begin
first_addr = 4'h1; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b10001001100: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10001001101: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b10001001110: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b10001001111: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b10001010000: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b10001010001: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b10001010010: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b10001010011: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b10001010100: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b10001010101: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b10001010110: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b10001010111: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b10001011000: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b10001011001: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b10001011010: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b10001011011: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b10001011100: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b10001011101: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b10001011110: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b10001011111: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b10001100000: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b10001100001: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b10001100010: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b10001100011: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b10001100100: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b10001100101: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b10001100110: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b10001100111: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b10001101000: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b10001101001: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b10001101010: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b10001101011: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b10001101100: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b10001101101: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b10001101110: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b10001101111: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b10001110000: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b10001110001: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b10001110010: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b10001110011: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b10001110100: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b10001110101: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b10001110110: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b10001110111: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b10001111000: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b10001111001: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b10001111010: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b10001111011: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b10001111100: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b10001111101: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b10001111110: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b10001111111: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b10010000000: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b10010000001: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b10010000010: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b10010000011: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b10010000100: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b10010000101: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b10010000110: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b10010000111: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b10010001000: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b10010001001: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b10010001010: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b10010001011: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b10010001100: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b10010001101: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b10010001110: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b10010001111: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b10010010000: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b10010010001: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b10010010010: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b10010010011: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b10010010100: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b10010010101: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b10010010110: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b10010010111: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b10010011000: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b10010011001: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b10010011010: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b10010011011: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b10010011100: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b10010011101: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b10010011110: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b10010011111: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b10010100000: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b10010100001: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b10010100010: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b10010100011: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b10010100100: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b10010100101: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b10010100110: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b10010100111: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b10010101000: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b10010101001: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b10010101010: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b10010101011: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b10010101100: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b10010101101: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b10010101110: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b10010101111: begin
first_addr = 4'h1; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b10010110000: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10010110001: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b10010110010: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b10010110011: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b10010110100: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b10010110101: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b10010110110: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b10010110111: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b10010111000: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b10010111001: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b10010111010: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b10010111011: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b10010111100: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b10010111101: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b10010111110: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b10010111111: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b10011000000: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b10011000001: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b10011000010: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b10011000011: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b10011000100: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b10011000101: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b10011000110: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b10011000111: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b10011001000: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b10011001001: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b10011001010: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b10011001011: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b10011001100: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b10011001101: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b10011001110: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b10011001111: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b10011010000: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b10011010001: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b10011010010: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b10011010011: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b10011010100: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b10011010101: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b10011010110: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b10011010111: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b10011011000: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b10011011001: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b10011011010: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b10011011011: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b10011011100: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b10011011101: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b10011011110: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b10011011111: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b10011100000: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b10011100001: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b10011100010: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b10011100011: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b10011100100: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b10011100101: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b10011100110: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b10011100111: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b10011101000: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b10011101001: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b10011101010: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b10011101011: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b10011101100: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b10011101101: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b10011101110: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b10011101111: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b10011110000: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b10011110001: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b10011110010: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b10011110011: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b10011110100: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b10011110101: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b10011110110: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b10011110111: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b10011111000: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b10011111001: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b10011111010: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b10011111011: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b10011111100: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b10011111101: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b10011111110: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b10011111111: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b10100000000: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b10100000001: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b10100000010: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b10100000011: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b10100000100: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b10100000101: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b10100000110: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b10100000111: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b10100001000: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b10100001001: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b10100001010: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b10100001011: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b10100001100: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b10100001101: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b10100001110: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b10100001111: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b10100010000: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b10100010001: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b10100010010: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b10100010011: begin
first_addr = 4'h1; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b10100010100: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10100010101: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b10100010110: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b10100010111: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b10100011000: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b10100011001: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b10100011010: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b10100011011: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b10100011100: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b10100011101: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b10100011110: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b10100011111: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b10100100000: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b10100100001: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b10100100010: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b10100100011: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b10100100100: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b10100100101: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b10100100110: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b10100100111: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b10100101000: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b10100101001: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b10100101010: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b10100101011: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b10100101100: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b10100101101: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b10100101110: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b10100101111: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b10100110000: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b10100110001: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b10100110010: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b10100110011: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b10100110100: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b10100110101: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b10100110110: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b10100110111: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b10100111000: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b10100111001: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b10100111010: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b10100111011: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b10100111100: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b10100111101: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b10100111110: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b10100111111: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b10101000000: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b10101000001: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b10101000010: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b10101000011: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b10101000100: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b10101000101: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b10101000110: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b10101000111: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b10101001000: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b10101001001: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b10101001010: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b10101001011: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b10101001100: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b10101001101: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b10101001110: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b10101001111: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b10101010000: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b10101010001: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b10101010010: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b10101010011: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b10101010100: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b10101010101: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b10101010110: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b10101010111: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b10101011000: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b10101011001: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b10101011010: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b10101011011: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b10101011100: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b10101011101: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b10101011110: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b10101011111: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b10101100000: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b10101100001: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b10101100010: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b10101100011: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b10101100100: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b10101100101: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b10101100110: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b10101100111: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b10101101000: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b10101101001: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b10101101010: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b10101101011: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b10101101100: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b10101101101: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b10101101110: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b10101101111: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b10101110000: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b10101110001: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b10101110010: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b10101110011: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b10101110100: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b10101110101: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b10101110110: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b10101110111: begin
first_addr = 4'h1; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b10101111000: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10101111001: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b10101111010: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b10101111011: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b10101111100: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b10101111101: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b10101111110: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b10101111111: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b10110000000: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b10110000001: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b10110000010: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b10110000011: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b10110000100: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b10110000101: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b10110000110: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b10110000111: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b10110001000: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b10110001001: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b10110001010: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b10110001011: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b10110001100: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b10110001101: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b10110001110: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b10110001111: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b10110010000: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b10110010001: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b10110010010: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b10110010011: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b10110010100: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b10110010101: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b10110010110: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b10110010111: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b10110011000: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b10110011001: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b10110011010: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b10110011011: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b10110011100: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b10110011101: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b10110011110: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b10110011111: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b10110100000: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b10110100001: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b10110100010: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b10110100011: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b10110100100: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b10110100101: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b10110100110: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b10110100111: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b10110101000: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b10110101001: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b10110101010: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b10110101011: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b10110101100: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b10110101101: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b10110101110: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b10110101111: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b10110110000: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b10110110001: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b10110110010: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b10110110011: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b10110110100: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b10110110101: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b10110110110: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b10110110111: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b10110111000: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b10110111001: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b10110111010: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b10110111011: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b10110111100: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b10110111101: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b10110111110: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b10110111111: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b10111000000: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b10111000001: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b10111000010: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b10111000011: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b10111000100: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b10111000101: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b10111000110: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b10111000111: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b10111001000: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b10111001001: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b10111001010: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b10111001011: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b10111001100: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b10111001101: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b10111001110: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b10111001111: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b10111010000: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b10111010001: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b10111010010: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b10111010011: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b10111010100: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b10111010101: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b10111010110: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b10111010111: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b10111011000: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b10111011001: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b10111011010: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b10111011011: begin
first_addr = 4'h1; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b10111011100: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b10111011101: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b10111011110: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b10111011111: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b10111100000: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b10111100001: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b10111100010: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b10111100011: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b10111100100: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b10111100101: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b10111100110: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b10111100111: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b10111101000: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b10111101001: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b10111101010: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b10111101011: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b10111101100: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b10111101101: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b10111101110: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b10111101111: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b10111110000: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b10111110001: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b10111110010: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b10111110011: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b10111110100: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b10111110101: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b10111110110: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b10111110111: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b10111111000: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b10111111001: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b10111111010: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b10111111011: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b10111111100: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b10111111101: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b10111111110: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b10111111111: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b11000000000: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b11000000001: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b11000000010: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b11000000011: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b11000000100: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b11000000101: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b11000000110: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b11000000111: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b11000001000: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b11000001001: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b11000001010: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b11000001011: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b11000001100: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b11000001101: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b11000001110: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b11000001111: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b11000010000: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b11000010001: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b11000010010: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b11000010011: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b11000010100: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b11000010101: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b11000010110: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b11000010111: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b11000011000: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b11000011001: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b11000011010: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b11000011011: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b11000011100: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b11000011101: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b11000011110: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b11000011111: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b11000100000: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b11000100001: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b11000100010: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b11000100011: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b11000100100: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b11000100101: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b11000100110: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b11000100111: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b11000101000: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b11000101001: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b11000101010: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b11000101011: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b11000101100: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b11000101101: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b11000101110: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b11000101111: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b11000110000: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b11000110001: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b11000110010: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b11000110011: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b11000110100: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b11000110101: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b11000110110: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b11000110111: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b11000111000: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b11000111001: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b11000111010: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b11000111011: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b11000111100: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b11000111101: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b11000111110: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b11000111111: begin
first_addr = 4'h1; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b11001000000: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11001000001: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b11001000010: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b11001000011: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b11001000100: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b11001000101: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b11001000110: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b11001000111: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b11001001000: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b11001001001: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b11001001010: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b11001001011: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b11001001100: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b11001001101: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b11001001110: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b11001001111: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b11001010000: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b11001010001: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b11001010010: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b11001010011: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b11001010100: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b11001010101: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b11001010110: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b11001010111: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b11001011000: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b11001011001: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b11001011010: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b11001011011: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b11001011100: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b11001011101: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b11001011110: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b11001011111: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b11001100000: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b11001100001: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b11001100010: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b11001100011: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b11001100100: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b11001100101: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b11001100110: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b11001100111: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b11001101000: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b11001101001: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b11001101010: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b11001101011: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b11001101100: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b11001101101: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b11001101110: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b11001101111: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b11001110000: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b11001110001: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b11001110010: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b11001110011: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b11001110100: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b11001110101: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b11001110110: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b11001110111: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b11001111000: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b11001111001: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b11001111010: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b11001111011: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b11001111100: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b11001111101: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b11001111110: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b11001111111: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b11010000000: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b11010000001: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b11010000010: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b11010000011: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b11010000100: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b11010000101: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b11010000110: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b11010000111: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b11010001000: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b11010001001: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b11010001010: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b11010001011: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b11010001100: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b11010001101: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b11010001110: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b11010001111: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b11010010000: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b11010010001: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b11010010010: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b11010010011: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b11010010100: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b11010010101: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b11010010110: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b11010010111: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b11010011000: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b11010011001: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b11010011010: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b11010011011: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b11010011100: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b11010011101: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b11010011110: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b11010011111: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b11010100000: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b11010100001: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b11010100010: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b11010100011: begin
first_addr = 4'h1; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b11010100100: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11010100101: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b11010100110: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b11010100111: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b11010101000: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b11010101001: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b11010101010: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b11010101011: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b11010101100: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b11010101101: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b11010101110: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b11010101111: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b11010110000: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b11010110001: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b11010110010: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b11010110011: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b11010110100: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b11010110101: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b11010110110: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b11010110111: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b11010111000: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b11010111001: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b11010111010: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b11010111011: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b11010111100: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b11010111101: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b11010111110: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b11010111111: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b11011000000: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b11011000001: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b11011000010: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b11011000011: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b11011000100: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b11011000101: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b11011000110: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b11011000111: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b11011001000: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b11011001001: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b11011001010: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b11011001011: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b11011001100: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b11011001101: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b11011001110: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b11011001111: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b11011010000: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b11011010001: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b11011010010: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b11011010011: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b11011010100: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b11011010101: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b11011010110: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b11011010111: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b11011011000: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b11011011001: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b11011011010: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b11011011011: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b11011011100: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b11011011101: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b11011011110: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b11011011111: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b11011100000: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b11011100001: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b11011100010: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b11011100011: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b11011100100: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b11011100101: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b11011100110: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b11011100111: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b11011101000: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b11011101001: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b11011101010: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b11011101011: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b11011101100: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b11011101101: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b11011101110: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b11011101111: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b11011110000: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b11011110001: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b11011110010: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b11011110011: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b11011110100: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b11011110101: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b11011110110: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b11011110111: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b11011111000: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b11011111001: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b11011111010: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b11011111011: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b11011111100: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b11011111101: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b11011111110: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b11011111111: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b11100000000: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b11100000001: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b11100000010: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b11100000011: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b11100000100: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b11100000101: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b11100000110: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b11100000111: begin
first_addr = 4'h1; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b11100001000: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11100001001: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b11100001010: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b11100001011: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b11100001100: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b11100001101: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b11100001110: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b11100001111: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b11100010000: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b11100010001: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b11100010010: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b11100010011: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b11100010100: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b11100010101: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b11100010110: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b11100010111: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b11100011000: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b11100011001: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b11100011010: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b11100011011: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b11100011100: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b11100011101: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b11100011110: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b11100011111: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b11100100000: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b11100100001: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b11100100010: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b11100100011: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b11100100100: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b11100100101: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b11100100110: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b11100100111: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b11100101000: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b11100101001: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b11100101010: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b11100101011: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b11100101100: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b11100101101: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b11100101110: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b11100101111: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b11100110000: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b11100110001: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b11100110010: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b11100110011: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b11100110100: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b11100110101: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b11100110110: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b11100110111: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b11100111000: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b11100111001: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b11100111010: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b11100111011: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b11100111100: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b11100111101: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b11100111110: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b11100111111: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b11101000000: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b11101000001: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b11101000010: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b11101000011: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b11101000100: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b11101000101: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b11101000110: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b11101000111: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b11101001000: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b11101001001: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b11101001010: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b11101001011: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b11101001100: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b11101001101: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b11101001110: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b11101001111: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b11101010000: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b11101010001: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b11101010010: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b11101010011: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b11101010100: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b11101010101: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b11101010110: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b11101010111: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b11101011000: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b11101011001: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b11101011010: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b11101011011: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b11101011100: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b11101011101: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b11101011110: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b11101011111: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b11101100000: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b11101100001: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b11101100010: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b11101100011: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b11101100100: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b11101100101: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b11101100110: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b11101100111: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b11101101000: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b11101101001: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b11101101010: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b11101101011: begin
first_addr = 4'h1; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b11101101100: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11101101101: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b11101101110: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b11101101111: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b11101110000: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b11101110001: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b11101110010: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b11101110011: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b11101110100: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b11101110101: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b11101110110: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b11101110111: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b11101111000: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b11101111001: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b11101111010: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b11101111011: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b11101111100: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b11101111101: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b11101111110: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b11101111111: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b11110000000: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b11110000001: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b11110000010: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b11110000011: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b11110000100: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b11110000101: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b11110000110: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b11110000111: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b11110001000: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b11110001001: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b11110001010: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b11110001011: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b11110001100: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b11110001101: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b11110001110: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b11110001111: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b11110010000: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b11110010001: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b11110010010: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b11110010011: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b11110010100: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b11110010101: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b11110010110: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b11110010111: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b11110011000: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b11110011001: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b11110011010: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b11110011011: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b11110011100: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b11110011101: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b11110011110: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b11110011111: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b11110100000: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b11110100001: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b11110100010: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b11110100011: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b11110100100: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b11110100101: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b11110100110: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b11110100111: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b11110101000: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b11110101001: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b11110101010: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b11110101011: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b11110101100: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b11110101101: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b11110101110: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b11110101111: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b11110110000: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b11110110001: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b11110110010: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b11110110011: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b11110110100: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b11110110101: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b11110110110: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b11110110111: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b11110111000: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b11110111001: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b11110111010: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b11110111011: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b11110111100: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b11110111101: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b11110111110: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b11110111111: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b11111000000: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b11111000001: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b11111000010: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b11111000011: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b11111000100: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b11111000101: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b11111000110: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b11111000111: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b11111001000: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b11111001001: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b11111001010: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b11111001011: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b11111001100: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b11111001101: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b11111001110: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b11111001111: begin
first_addr = 4'h1; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b11111010000: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b11111010001: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b11111010010: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b11111010011: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b11111010100: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b11111010101: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b11111010110: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b11111010111: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b11111011000: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b11111011001: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b11111011010: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b11111011011: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b11111011100: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b11111011101: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b11111011110: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b11111011111: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b11111100000: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b11111100001: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b11111100010: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b11111100011: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b11111100100: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b11111100101: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b11111100110: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b11111100111: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b11111101000: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b11111101001: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b11111101010: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b11111101011: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b11111101100: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b11111101101: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b11111101110: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b11111101111: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b11111110000: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b11111110001: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b11111110010: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b11111110011: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b11111110100: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b11111110101: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b11111110110: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b11111110111: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b11111111000: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b11111111001: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b11111111010: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b11111111011: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b11111111100: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b11111111101: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b11111111110: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b11111111111: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b100000000000: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b100000000001: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b100000000010: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b100000000011: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b100000000100: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b100000000101: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b100000000110: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b100000000111: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b100000001000: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b100000001001: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b100000001010: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b100000001011: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b100000001100: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b100000001101: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b100000001110: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b100000001111: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b100000010000: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b100000010001: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b100000010010: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b100000010011: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b100000010100: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b100000010101: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b100000010110: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b100000010111: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b100000011000: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b100000011001: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b100000011010: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b100000011011: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b100000011100: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b100000011101: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b100000011110: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b100000011111: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b100000100000: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b100000100001: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b100000100010: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b100000100011: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b100000100100: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b100000100101: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b100000100110: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b100000100111: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b100000101000: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b100000101001: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b100000101010: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b100000101011: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b100000101100: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b100000101101: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b100000101110: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b100000101111: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b100000110000: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b100000110001: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b100000110010: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b100000110011: begin
first_addr = 4'h2; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b100000110100: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100000110101: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b100000110110: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b100000110111: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b100000111000: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b100000111001: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b100000111010: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b100000111011: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b100000111100: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b100000111101: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b100000111110: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b100000111111: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b100001000000: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b100001000001: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b100001000010: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b100001000011: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b100001000100: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b100001000101: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b100001000110: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b100001000111: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b100001001000: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b100001001001: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b100001001010: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b100001001011: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b100001001100: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b100001001101: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b100001001110: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b100001001111: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b100001010000: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b100001010001: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b100001010010: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b100001010011: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b100001010100: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b100001010101: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b100001010110: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b100001010111: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b100001011000: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b100001011001: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b100001011010: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b100001011011: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b100001011100: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b100001011101: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b100001011110: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b100001011111: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b100001100000: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b100001100001: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b100001100010: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b100001100011: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b100001100100: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b100001100101: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b100001100110: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b100001100111: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b100001101000: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b100001101001: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b100001101010: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b100001101011: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b100001101100: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b100001101101: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b100001101110: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b100001101111: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b100001110000: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b100001110001: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b100001110010: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b100001110011: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b100001110100: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b100001110101: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b100001110110: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b100001110111: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b100001111000: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b100001111001: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b100001111010: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b100001111011: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b100001111100: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b100001111101: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b100001111110: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b100001111111: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b100010000000: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b100010000001: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b100010000010: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b100010000011: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b100010000100: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b100010000101: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b100010000110: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b100010000111: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b100010001000: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b100010001001: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b100010001010: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b100010001011: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b100010001100: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b100010001101: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b100010001110: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b100010001111: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b100010010000: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b100010010001: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b100010010010: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b100010010011: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b100010010100: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b100010010101: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b100010010110: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b100010010111: begin
first_addr = 4'h2; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b100010011000: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100010011001: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b100010011010: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b100010011011: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b100010011100: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b100010011101: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b100010011110: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b100010011111: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b100010100000: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b100010100001: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b100010100010: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b100010100011: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b100010100100: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b100010100101: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b100010100110: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b100010100111: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b100010101000: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b100010101001: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b100010101010: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b100010101011: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b100010101100: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b100010101101: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b100010101110: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b100010101111: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b100010110000: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b100010110001: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b100010110010: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b100010110011: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b100010110100: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b100010110101: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b100010110110: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b100010110111: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b100010111000: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b100010111001: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b100010111010: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b100010111011: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b100010111100: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b100010111101: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b100010111110: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b100010111111: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b100011000000: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b100011000001: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b100011000010: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b100011000011: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b100011000100: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b100011000101: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b100011000110: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b100011000111: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b100011001000: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b100011001001: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b100011001010: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b100011001011: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b100011001100: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b100011001101: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b100011001110: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b100011001111: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b100011010000: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b100011010001: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b100011010010: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b100011010011: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b100011010100: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b100011010101: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b100011010110: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b100011010111: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b100011011000: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b100011011001: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b100011011010: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b100011011011: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b100011011100: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b100011011101: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b100011011110: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b100011011111: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b100011100000: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b100011100001: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b100011100010: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b100011100011: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b100011100100: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b100011100101: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b100011100110: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b100011100111: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b100011101000: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b100011101001: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b100011101010: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b100011101011: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b100011101100: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b100011101101: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b100011101110: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b100011101111: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b100011110000: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b100011110001: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b100011110010: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b100011110011: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b100011110100: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b100011110101: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b100011110110: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b100011110111: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b100011111000: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b100011111001: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b100011111010: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b100011111011: begin
first_addr = 4'h2; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b100011111100: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100011111101: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b100011111110: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b100011111111: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b100100000000: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b100100000001: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b100100000010: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b100100000011: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b100100000100: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b100100000101: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b100100000110: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b100100000111: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b100100001000: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b100100001001: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b100100001010: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b100100001011: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b100100001100: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b100100001101: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b100100001110: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b100100001111: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b100100010000: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b100100010001: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b100100010010: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b100100010011: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b100100010100: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b100100010101: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b100100010110: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b100100010111: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b100100011000: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b100100011001: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b100100011010: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b100100011011: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b100100011100: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b100100011101: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b100100011110: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b100100011111: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b100100100000: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b100100100001: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b100100100010: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b100100100011: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b100100100100: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b100100100101: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b100100100110: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b100100100111: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b100100101000: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b100100101001: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b100100101010: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b100100101011: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b100100101100: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b100100101101: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b100100101110: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b100100101111: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b100100110000: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b100100110001: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b100100110010: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b100100110011: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b100100110100: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b100100110101: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b100100110110: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b100100110111: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b100100111000: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b100100111001: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b100100111010: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b100100111011: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b100100111100: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b100100111101: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b100100111110: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b100100111111: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b100101000000: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b100101000001: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b100101000010: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b100101000011: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b100101000100: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b100101000101: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b100101000110: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b100101000111: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b100101001000: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b100101001001: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b100101001010: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b100101001011: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b100101001100: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b100101001101: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b100101001110: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b100101001111: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b100101010000: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b100101010001: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b100101010010: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b100101010011: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b100101010100: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b100101010101: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b100101010110: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b100101010111: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b100101011000: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b100101011001: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b100101011010: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b100101011011: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b100101011100: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b100101011101: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b100101011110: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b100101011111: begin
first_addr = 4'h2; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b100101100000: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100101100001: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b100101100010: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b100101100011: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b100101100100: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b100101100101: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b100101100110: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b100101100111: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b100101101000: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b100101101001: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b100101101010: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b100101101011: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b100101101100: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b100101101101: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b100101101110: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b100101101111: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b100101110000: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b100101110001: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b100101110010: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b100101110011: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b100101110100: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b100101110101: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b100101110110: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b100101110111: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b100101111000: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b100101111001: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b100101111010: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b100101111011: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b100101111100: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b100101111101: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b100101111110: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b100101111111: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b100110000000: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b100110000001: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b100110000010: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b100110000011: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b100110000100: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b100110000101: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b100110000110: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b100110000111: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b100110001000: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b100110001001: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b100110001010: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b100110001011: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b100110001100: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b100110001101: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b100110001110: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b100110001111: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b100110010000: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b100110010001: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b100110010010: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b100110010011: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b100110010100: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b100110010101: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b100110010110: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b100110010111: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b100110011000: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b100110011001: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b100110011010: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b100110011011: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b100110011100: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b100110011101: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b100110011110: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b100110011111: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b100110100000: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b100110100001: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b100110100010: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b100110100011: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b100110100100: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b100110100101: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b100110100110: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b100110100111: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b100110101000: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b100110101001: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b100110101010: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b100110101011: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b100110101100: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b100110101101: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b100110101110: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b100110101111: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b100110110000: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b100110110001: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b100110110010: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b100110110011: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b100110110100: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b100110110101: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b100110110110: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b100110110111: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b100110111000: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b100110111001: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b100110111010: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b100110111011: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b100110111100: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b100110111101: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b100110111110: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b100110111111: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b100111000000: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b100111000001: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b100111000010: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b100111000011: begin
first_addr = 4'h2; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b100111000100: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b100111000101: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b100111000110: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b100111000111: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b100111001000: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b100111001001: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b100111001010: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b100111001011: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b100111001100: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b100111001101: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b100111001110: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b100111001111: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b100111010000: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b100111010001: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b100111010010: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b100111010011: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b100111010100: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b100111010101: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b100111010110: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b100111010111: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b100111011000: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b100111011001: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b100111011010: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b100111011011: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b100111011100: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b100111011101: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b100111011110: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b100111011111: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b100111100000: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b100111100001: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b100111100010: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b100111100011: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b100111100100: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b100111100101: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b100111100110: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b100111100111: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b100111101000: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b100111101001: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b100111101010: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b100111101011: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b100111101100: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b100111101101: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b100111101110: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b100111101111: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b100111110000: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b100111110001: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b100111110010: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b100111110011: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b100111110100: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b100111110101: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b100111110110: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b100111110111: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b100111111000: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b100111111001: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b100111111010: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b100111111011: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b100111111100: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b100111111101: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b100111111110: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b100111111111: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b101000000000: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b101000000001: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b101000000010: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b101000000011: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b101000000100: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b101000000101: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b101000000110: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b101000000111: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b101000001000: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b101000001001: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b101000001010: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b101000001011: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b101000001100: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b101000001101: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b101000001110: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b101000001111: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b101000010000: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b101000010001: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b101000010010: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b101000010011: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b101000010100: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b101000010101: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b101000010110: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b101000010111: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b101000011000: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b101000011001: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b101000011010: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b101000011011: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b101000011100: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b101000011101: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b101000011110: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b101000011111: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b101000100000: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b101000100001: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b101000100010: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b101000100011: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b101000100100: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b101000100101: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b101000100110: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b101000100111: begin
first_addr = 4'h2; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b101000101000: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101000101001: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b101000101010: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b101000101011: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b101000101100: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b101000101101: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b101000101110: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b101000101111: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b101000110000: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b101000110001: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b101000110010: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b101000110011: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b101000110100: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b101000110101: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b101000110110: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b101000110111: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b101000111000: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b101000111001: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b101000111010: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b101000111011: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b101000111100: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b101000111101: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b101000111110: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b101000111111: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b101001000000: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b101001000001: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b101001000010: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b101001000011: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b101001000100: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b101001000101: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b101001000110: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b101001000111: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b101001001000: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b101001001001: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b101001001010: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b101001001011: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b101001001100: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b101001001101: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b101001001110: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b101001001111: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b101001010000: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b101001010001: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b101001010010: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b101001010011: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b101001010100: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b101001010101: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b101001010110: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b101001010111: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b101001011000: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b101001011001: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b101001011010: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b101001011011: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b101001011100: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b101001011101: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b101001011110: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b101001011111: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b101001100000: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b101001100001: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b101001100010: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b101001100011: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b101001100100: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b101001100101: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b101001100110: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b101001100111: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b101001101000: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b101001101001: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b101001101010: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b101001101011: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b101001101100: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b101001101101: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b101001101110: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b101001101111: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b101001110000: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b101001110001: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b101001110010: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b101001110011: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b101001110100: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b101001110101: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b101001110110: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b101001110111: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b101001111000: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b101001111001: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b101001111010: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b101001111011: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b101001111100: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b101001111101: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b101001111110: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b101001111111: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b101010000000: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b101010000001: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b101010000010: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b101010000011: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b101010000100: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b101010000101: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b101010000110: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b101010000111: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b101010001000: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b101010001001: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b101010001010: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b101010001011: begin
first_addr = 4'h2; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b101010001100: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101010001101: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b101010001110: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b101010001111: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b101010010000: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b101010010001: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b101010010010: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b101010010011: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b101010010100: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b101010010101: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b101010010110: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b101010010111: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b101010011000: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b101010011001: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b101010011010: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b101010011011: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b101010011100: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b101010011101: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b101010011110: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b101010011111: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b101010100000: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b101010100001: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b101010100010: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b101010100011: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b101010100100: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b101010100101: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b101010100110: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b101010100111: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b101010101000: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b101010101001: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b101010101010: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b101010101011: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b101010101100: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b101010101101: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b101010101110: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b101010101111: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b101010110000: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b101010110001: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b101010110010: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b101010110011: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b101010110100: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b101010110101: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b101010110110: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b101010110111: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b101010111000: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b101010111001: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b101010111010: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b101010111011: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b101010111100: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b101010111101: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b101010111110: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b101010111111: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b101011000000: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b101011000001: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b101011000010: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b101011000011: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b101011000100: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b101011000101: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b101011000110: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b101011000111: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b101011001000: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b101011001001: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b101011001010: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b101011001011: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b101011001100: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b101011001101: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b101011001110: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b101011001111: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b101011010000: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b101011010001: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b101011010010: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b101011010011: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b101011010100: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b101011010101: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b101011010110: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b101011010111: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b101011011000: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b101011011001: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b101011011010: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b101011011011: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b101011011100: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b101011011101: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b101011011110: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b101011011111: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b101011100000: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b101011100001: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b101011100010: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b101011100011: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b101011100100: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b101011100101: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b101011100110: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b101011100111: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b101011101000: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b101011101001: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b101011101010: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b101011101011: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b101011101100: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b101011101101: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b101011101110: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b101011101111: begin
first_addr = 4'h2; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b101011110000: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101011110001: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b101011110010: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b101011110011: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b101011110100: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b101011110101: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b101011110110: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b101011110111: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b101011111000: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b101011111001: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b101011111010: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b101011111011: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b101011111100: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b101011111101: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b101011111110: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b101011111111: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b101100000000: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b101100000001: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b101100000010: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b101100000011: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b101100000100: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b101100000101: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b101100000110: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b101100000111: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b101100001000: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b101100001001: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b101100001010: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b101100001011: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b101100001100: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b101100001101: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b101100001110: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b101100001111: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b101100010000: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b101100010001: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b101100010010: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b101100010011: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b101100010100: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b101100010101: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b101100010110: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b101100010111: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b101100011000: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b101100011001: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b101100011010: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b101100011011: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b101100011100: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b101100011101: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b101100011110: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b101100011111: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b101100100000: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b101100100001: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b101100100010: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b101100100011: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b101100100100: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b101100100101: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b101100100110: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b101100100111: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b101100101000: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b101100101001: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b101100101010: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b101100101011: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b101100101100: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b101100101101: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b101100101110: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b101100101111: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b101100110000: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b101100110001: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b101100110010: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b101100110011: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b101100110100: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b101100110101: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b101100110110: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b101100110111: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b101100111000: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b101100111001: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b101100111010: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b101100111011: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b101100111100: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b101100111101: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b101100111110: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b101100111111: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b101101000000: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b101101000001: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b101101000010: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b101101000011: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b101101000100: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b101101000101: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b101101000110: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b101101000111: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b101101001000: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b101101001001: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b101101001010: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b101101001011: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b101101001100: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b101101001101: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b101101001110: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b101101001111: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b101101010000: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b101101010001: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b101101010010: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b101101010011: begin
first_addr = 4'h2; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b101101010100: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101101010101: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b101101010110: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b101101010111: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b101101011000: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b101101011001: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b101101011010: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b101101011011: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b101101011100: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b101101011101: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b101101011110: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b101101011111: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b101101100000: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b101101100001: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b101101100010: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b101101100011: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b101101100100: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b101101100101: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b101101100110: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b101101100111: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b101101101000: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b101101101001: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b101101101010: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b101101101011: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b101101101100: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b101101101101: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b101101101110: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b101101101111: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b101101110000: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b101101110001: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b101101110010: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b101101110011: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b101101110100: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b101101110101: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b101101110110: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b101101110111: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b101101111000: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b101101111001: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b101101111010: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b101101111011: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b101101111100: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b101101111101: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b101101111110: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b101101111111: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b101110000000: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b101110000001: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b101110000010: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b101110000011: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b101110000100: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b101110000101: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b101110000110: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b101110000111: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b101110001000: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b101110001001: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b101110001010: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b101110001011: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b101110001100: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b101110001101: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b101110001110: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b101110001111: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b101110010000: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b101110010001: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b101110010010: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b101110010011: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b101110010100: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b101110010101: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b101110010110: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b101110010111: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b101110011000: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b101110011001: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b101110011010: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b101110011011: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b101110011100: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b101110011101: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b101110011110: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b101110011111: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b101110100000: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b101110100001: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b101110100010: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b101110100011: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b101110100100: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b101110100101: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b101110100110: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b101110100111: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b101110101000: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b101110101001: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b101110101010: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b101110101011: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b101110101100: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b101110101101: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b101110101110: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b101110101111: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b101110110000: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b101110110001: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b101110110010: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b101110110011: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b101110110100: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b101110110101: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b101110110110: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b101110110111: begin
first_addr = 4'h2; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b101110111000: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b101110111001: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b101110111010: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b101110111011: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b101110111100: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b101110111101: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b101110111110: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b101110111111: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b101111000000: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b101111000001: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b101111000010: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b101111000011: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b101111000100: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b101111000101: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b101111000110: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b101111000111: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b101111001000: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b101111001001: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b101111001010: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b101111001011: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b101111001100: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b101111001101: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b101111001110: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b101111001111: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b101111010000: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b101111010001: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b101111010010: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b101111010011: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b101111010100: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b101111010101: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b101111010110: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b101111010111: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b101111011000: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b101111011001: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b101111011010: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b101111011011: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b101111011100: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b101111011101: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b101111011110: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b101111011111: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b101111100000: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b101111100001: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b101111100010: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b101111100011: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b101111100100: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b101111100101: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b101111100110: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b101111100111: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b101111101000: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b101111101001: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b101111101010: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b101111101011: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b101111101100: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b101111101101: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b101111101110: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b101111101111: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b101111110000: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b101111110001: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b101111110010: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b101111110011: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b101111110100: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b101111110101: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b101111110110: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b101111110111: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b101111111000: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b101111111001: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b101111111010: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b101111111011: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b101111111100: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b101111111101: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b101111111110: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b101111111111: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b110000000000: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b110000000001: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b110000000010: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b110000000011: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b110000000100: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b110000000101: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b110000000110: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b110000000111: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b110000001000: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b110000001001: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b110000001010: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b110000001011: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b110000001100: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b110000001101: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b110000001110: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b110000001111: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b110000010000: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b110000010001: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b110000010010: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b110000010011: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b110000010100: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b110000010101: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b110000010110: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b110000010111: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b110000011000: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b110000011001: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b110000011010: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b110000011011: begin
first_addr = 4'h3; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b110000011100: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110000011101: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b110000011110: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b110000011111: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b110000100000: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b110000100001: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b110000100010: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b110000100011: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b110000100100: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b110000100101: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b110000100110: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b110000100111: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b110000101000: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b110000101001: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b110000101010: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b110000101011: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b110000101100: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b110000101101: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b110000101110: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b110000101111: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b110000110000: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b110000110001: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b110000110010: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b110000110011: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b110000110100: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b110000110101: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b110000110110: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b110000110111: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b110000111000: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b110000111001: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b110000111010: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b110000111011: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b110000111100: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b110000111101: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b110000111110: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b110000111111: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b110001000000: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b110001000001: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b110001000010: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b110001000011: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b110001000100: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b110001000101: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b110001000110: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b110001000111: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b110001001000: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b110001001001: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b110001001010: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b110001001011: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b110001001100: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b110001001101: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b110001001110: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b110001001111: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b110001010000: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b110001010001: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b110001010010: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b110001010011: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b110001010100: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b110001010101: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b110001010110: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b110001010111: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b110001011000: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b110001011001: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b110001011010: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b110001011011: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b110001011100: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b110001011101: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b110001011110: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b110001011111: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b110001100000: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b110001100001: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b110001100010: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b110001100011: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b110001100100: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b110001100101: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b110001100110: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b110001100111: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b110001101000: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b110001101001: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b110001101010: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b110001101011: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b110001101100: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b110001101101: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b110001101110: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b110001101111: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b110001110000: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b110001110001: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b110001110010: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b110001110011: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b110001110100: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b110001110101: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b110001110110: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b110001110111: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b110001111000: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b110001111001: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b110001111010: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b110001111011: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b110001111100: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b110001111101: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b110001111110: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b110001111111: begin
first_addr = 4'h3; 
second_addr = 4'h1; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b110010000000: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110010000001: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b110010000010: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b110010000011: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b110010000100: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b110010000101: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b110010000110: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b110010000111: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b110010001000: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b110010001001: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b110010001010: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b110010001011: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b110010001100: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b110010001101: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b110010001110: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b110010001111: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b110010010000: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b110010010001: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b110010010010: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b110010010011: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b110010010100: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b110010010101: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b110010010110: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b110010010111: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b110010011000: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b110010011001: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b110010011010: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b110010011011: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b110010011100: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b110010011101: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b110010011110: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b110010011111: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b110010100000: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b110010100001: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b110010100010: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b110010100011: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b110010100100: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b110010100101: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b110010100110: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b110010100111: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b110010101000: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b110010101001: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b110010101010: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b110010101011: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b110010101100: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b110010101101: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b110010101110: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b110010101111: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b110010110000: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b110010110001: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b110010110010: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b110010110011: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b110010110100: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b110010110101: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b110010110110: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b110010110111: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b110010111000: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b110010111001: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b110010111010: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b110010111011: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b110010111100: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b110010111101: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b110010111110: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b110010111111: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b110011000000: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b110011000001: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b110011000010: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b110011000011: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b110011000100: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b110011000101: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b110011000110: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b110011000111: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b110011001000: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b110011001001: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b110011001010: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b110011001011: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b110011001100: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b110011001101: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b110011001110: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b110011001111: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b110011010000: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b110011010001: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b110011010010: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b110011010011: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b110011010100: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b110011010101: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b110011010110: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b110011010111: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b110011011000: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b110011011001: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b110011011010: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b110011011011: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b110011011100: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b110011011101: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b110011011110: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b110011011111: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b110011100000: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b110011100001: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b110011100010: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b110011100011: begin
first_addr = 4'h3; 
second_addr = 4'h2; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b110011100100: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110011100101: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b110011100110: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b110011100111: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b110011101000: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b110011101001: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b110011101010: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b110011101011: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b110011101100: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b110011101101: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b110011101110: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b110011101111: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b110011110000: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b110011110001: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b110011110010: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b110011110011: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b110011110100: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b110011110101: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b110011110110: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b110011110111: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b110011111000: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b110011111001: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b110011111010: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b110011111011: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b110011111100: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b110011111101: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b110011111110: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b110011111111: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b110100000000: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b110100000001: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b110100000010: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b110100000011: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b110100000100: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b110100000101: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b110100000110: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b110100000111: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b110100001000: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b110100001001: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b110100001010: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b110100001011: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b110100001100: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b110100001101: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b110100001110: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b110100001111: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b110100010000: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b110100010001: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b110100010010: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b110100010011: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b110100010100: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b110100010101: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b110100010110: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b110100010111: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b110100011000: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b110100011001: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b110100011010: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b110100011011: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b110100011100: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b110100011101: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b110100011110: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b110100011111: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b110100100000: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b110100100001: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b110100100010: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b110100100011: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b110100100100: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b110100100101: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b110100100110: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b110100100111: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b110100101000: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b110100101001: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b110100101010: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b110100101011: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b110100101100: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b110100101101: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b110100101110: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b110100101111: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b110100110000: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b110100110001: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b110100110010: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b110100110011: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b110100110100: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b110100110101: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b110100110110: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b110100110111: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b110100111000: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b110100111001: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b110100111010: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b110100111011: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b110100111100: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b110100111101: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b110100111110: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b110100111111: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b110101000000: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b110101000001: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b110101000010: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b110101000011: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b110101000100: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b110101000101: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b110101000110: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b110101000111: begin
first_addr = 4'h3; 
second_addr = 4'h3; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b110101001000: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110101001001: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b110101001010: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b110101001011: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b110101001100: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b110101001101: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b110101001110: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b110101001111: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b110101010000: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b110101010001: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b110101010010: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b110101010011: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b110101010100: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b110101010101: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b110101010110: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b110101010111: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b110101011000: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b110101011001: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b110101011010: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b110101011011: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b110101011100: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b110101011101: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b110101011110: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b110101011111: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b110101100000: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b110101100001: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b110101100010: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b110101100011: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b110101100100: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b110101100101: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b110101100110: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b110101100111: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b110101101000: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b110101101001: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b110101101010: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b110101101011: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b110101101100: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b110101101101: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b110101101110: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b110101101111: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b110101110000: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b110101110001: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b110101110010: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b110101110011: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b110101110100: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b110101110101: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b110101110110: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b110101110111: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b110101111000: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b110101111001: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b110101111010: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b110101111011: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b110101111100: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b110101111101: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b110101111110: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b110101111111: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b110110000000: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b110110000001: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b110110000010: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b110110000011: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b110110000100: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b110110000101: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b110110000110: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b110110000111: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b110110001000: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b110110001001: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b110110001010: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b110110001011: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b110110001100: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b110110001101: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b110110001110: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b110110001111: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b110110010000: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b110110010001: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b110110010010: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b110110010011: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b110110010100: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b110110010101: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b110110010110: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b110110010111: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b110110011000: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b110110011001: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b110110011010: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b110110011011: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b110110011100: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b110110011101: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b110110011110: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b110110011111: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b110110100000: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b110110100001: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b110110100010: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b110110100011: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b110110100100: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b110110100101: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b110110100110: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b110110100111: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b110110101000: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b110110101001: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b110110101010: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b110110101011: begin
first_addr = 4'h3; 
second_addr = 4'h4; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b110110101100: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b110110101101: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b110110101110: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b110110101111: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b110110110000: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b110110110001: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b110110110010: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b110110110011: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b110110110100: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b110110110101: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b110110110110: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b110110110111: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b110110111000: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b110110111001: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b110110111010: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b110110111011: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b110110111100: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b110110111101: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b110110111110: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b110110111111: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b110111000000: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b110111000001: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b110111000010: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b110111000011: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b110111000100: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b110111000101: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b110111000110: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b110111000111: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b110111001000: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b110111001001: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b110111001010: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b110111001011: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b110111001100: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b110111001101: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b110111001110: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b110111001111: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b110111010000: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b110111010001: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b110111010010: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b110111010011: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b110111010100: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b110111010101: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b110111010110: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b110111010111: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b110111011000: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b110111011001: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b110111011010: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b110111011011: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b110111011100: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b110111011101: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b110111011110: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b110111011111: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b110111100000: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b110111100001: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b110111100010: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b110111100011: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b110111100100: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b110111100101: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b110111100110: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b110111100111: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b110111101000: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b110111101001: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b110111101010: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b110111101011: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b110111101100: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b110111101101: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b110111101110: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b110111101111: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b110111110000: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b110111110001: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b110111110010: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b110111110011: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b110111110100: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b110111110101: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b110111110110: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b110111110111: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b110111111000: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b110111111001: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b110111111010: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b110111111011: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b110111111100: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b110111111101: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b110111111110: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b110111111111: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b111000000000: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b111000000001: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b111000000010: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b111000000011: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b111000000100: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b111000000101: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b111000000110: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b111000000111: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b111000001000: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b111000001001: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b111000001010: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b111000001011: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b111000001100: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b111000001101: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b111000001110: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b111000001111: begin
first_addr = 4'h3; 
second_addr = 4'h5; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b111000010000: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111000010001: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b111000010010: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b111000010011: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b111000010100: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b111000010101: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b111000010110: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b111000010111: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b111000011000: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b111000011001: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b111000011010: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b111000011011: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b111000011100: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b111000011101: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b111000011110: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b111000011111: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b111000100000: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b111000100001: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b111000100010: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b111000100011: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b111000100100: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b111000100101: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b111000100110: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b111000100111: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b111000101000: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b111000101001: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b111000101010: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b111000101011: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b111000101100: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b111000101101: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b111000101110: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b111000101111: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b111000110000: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b111000110001: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b111000110010: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b111000110011: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b111000110100: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b111000110101: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b111000110110: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b111000110111: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b111000111000: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b111000111001: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b111000111010: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b111000111011: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b111000111100: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b111000111101: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b111000111110: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b111000111111: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b111001000000: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b111001000001: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b111001000010: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b111001000011: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b111001000100: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b111001000101: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b111001000110: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b111001000111: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b111001001000: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b111001001001: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b111001001010: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b111001001011: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b111001001100: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b111001001101: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b111001001110: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b111001001111: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b111001010000: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b111001010001: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b111001010010: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b111001010011: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b111001010100: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b111001010101: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b111001010110: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b111001010111: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b111001011000: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b111001011001: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b111001011010: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b111001011011: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b111001011100: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b111001011101: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b111001011110: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b111001011111: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b111001100000: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b111001100001: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b111001100010: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b111001100011: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b111001100100: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b111001100101: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b111001100110: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b111001100111: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b111001101000: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b111001101001: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b111001101010: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b111001101011: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b111001101100: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b111001101101: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b111001101110: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b111001101111: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b111001110000: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b111001110001: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b111001110010: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b111001110011: begin
first_addr = 4'h3; 
second_addr = 4'h6; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b111001110100: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111001110101: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b111001110110: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b111001110111: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b111001111000: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b111001111001: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b111001111010: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b111001111011: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b111001111100: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b111001111101: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b111001111110: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b111001111111: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b111010000000: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b111010000001: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b111010000010: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b111010000011: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b111010000100: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b111010000101: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b111010000110: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b111010000111: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b111010001000: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b111010001001: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b111010001010: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b111010001011: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b111010001100: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b111010001101: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b111010001110: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b111010001111: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b111010010000: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b111010010001: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b111010010010: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b111010010011: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b111010010100: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b111010010101: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b111010010110: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b111010010111: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b111010011000: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b111010011001: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b111010011010: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b111010011011: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b111010011100: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b111010011101: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b111010011110: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b111010011111: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b111010100000: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b111010100001: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b111010100010: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b111010100011: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b111010100100: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b111010100101: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b111010100110: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b111010100111: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b111010101000: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b111010101001: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b111010101010: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b111010101011: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b111010101100: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b111010101101: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b111010101110: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b111010101111: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b111010110000: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b111010110001: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b111010110010: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b111010110011: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b111010110100: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b111010110101: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b111010110110: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b111010110111: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b111010111000: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b111010111001: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b111010111010: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b111010111011: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b111010111100: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b111010111101: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b111010111110: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b111010111111: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b111011000000: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b111011000001: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b111011000010: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b111011000011: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b111011000100: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b111011000101: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b111011000110: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b111011000111: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b111011001000: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b111011001001: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b111011001010: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b111011001011: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b111011001100: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b111011001101: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b111011001110: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b111011001111: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b111011010000: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b111011010001: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b111011010010: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b111011010011: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b111011010100: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b111011010101: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b111011010110: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b111011010111: begin
first_addr = 4'h3; 
second_addr = 4'h7; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b111011011000: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111011011001: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b111011011010: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b111011011011: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b111011011100: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b111011011101: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b111011011110: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b111011011111: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b111011100000: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b111011100001: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b111011100010: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b111011100011: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b111011100100: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b111011100101: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b111011100110: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b111011100111: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b111011101000: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b111011101001: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b111011101010: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b111011101011: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b111011101100: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b111011101101: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b111011101110: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b111011101111: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b111011110000: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b111011110001: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b111011110010: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b111011110011: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b111011110100: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b111011110101: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b111011110110: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b111011110111: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b111011111000: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b111011111001: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b111011111010: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b111011111011: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b111011111100: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b111011111101: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b111011111110: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b111011111111: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b111100000000: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b111100000001: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b111100000010: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b111100000011: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b111100000100: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b111100000101: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b111100000110: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b111100000111: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b111100001000: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b111100001001: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b111100001010: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b111100001011: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b111100001100: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b111100001101: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b111100001110: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b111100001111: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b111100010000: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b111100010001: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b111100010010: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b111100010011: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b111100010100: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b111100010101: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b111100010110: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b111100010111: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b111100011000: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b111100011001: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b111100011010: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b111100011011: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b111100011100: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b111100011101: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b111100011110: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b111100011111: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b111100100000: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b111100100001: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b111100100010: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b111100100011: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b111100100100: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b111100100101: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b111100100110: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b111100100111: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b111100101000: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b111100101001: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b111100101010: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b111100101011: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b111100101100: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b111100101101: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b111100101110: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b111100101111: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b111100110000: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b111100110001: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b111100110010: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b111100110011: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b111100110100: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b111100110101: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b111100110110: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b111100110111: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b111100111000: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b111100111001: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b111100111010: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b111100111011: begin
first_addr = 4'h3; 
second_addr = 4'h8; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b111100111100: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111100111101: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b111100111110: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b111100111111: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b111101000000: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b111101000001: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b111101000010: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b111101000011: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b111101000100: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b111101000101: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b111101000110: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b111101000111: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b111101001000: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b111101001001: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b111101001010: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b111101001011: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b111101001100: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b111101001101: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b111101001110: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b111101001111: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b111101010000: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b111101010001: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b111101010010: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b111101010011: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b111101010100: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b111101010101: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b111101010110: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b111101010111: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b111101011000: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b111101011001: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b111101011010: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b111101011011: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b111101011100: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b111101011101: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b111101011110: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b111101011111: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b111101100000: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b111101100001: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b111101100010: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b111101100011: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b111101100100: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b111101100101: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b111101100110: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b111101100111: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b111101101000: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b111101101001: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b111101101010: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b111101101011: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b111101101100: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b111101101101: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b111101101110: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b111101101111: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b111101110000: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b111101110001: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b111101110010: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b111101110011: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b111101110100: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b111101110101: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b111101110110: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b111101110111: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b111101111000: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b111101111001: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b111101111010: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b111101111011: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b111101111100: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b111101111101: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b111101111110: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b111101111111: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b111110000000: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b111110000001: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b111110000010: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b111110000011: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b111110000100: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b111110000101: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b111110000110: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b111110000111: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b111110001000: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b111110001001: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b111110001010: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b111110001011: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b111110001100: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b111110001101: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b111110001110: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b111110001111: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b111110010000: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b111110010001: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b111110010010: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b111110010011: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b111110010100: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b111110010101: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b111110010110: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b111110010111: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b111110011000: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b111110011001: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b111110011010: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b111110011011: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end

 10'b111110011100: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h6; 
end

 10'b111110011101: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h7; 
end

 10'b111110011110: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h8; 
end

 10'b111110011111: begin
first_addr = 4'h3; 
second_addr = 4'h9; 
third_addr = 4'h9; 
fourth_addr =4'h9; 
end

 10'b111110100000: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h0; 
end

 10'b111110100001: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h1; 
end

 10'b111110100010: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h2; 
end

 10'b111110100011: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h3; 
end

 10'b111110100100: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h4; 
end

 10'b111110100101: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h5; 
end

 10'b111110100110: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h6; 
end

 10'b111110100111: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h7; 
end

 10'b111110101000: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h8; 
end

 10'b111110101001: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h0; 
fourth_addr =4'h9; 
end

 10'b111110101010: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h0; 
end

 10'b111110101011: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h1; 
end

 10'b111110101100: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h2; 
end

 10'b111110101101: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h3; 
end

 10'b111110101110: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h4; 
end

 10'b111110101111: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h5; 
end

 10'b111110110000: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h6; 
end

 10'b111110110001: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h7; 
end

 10'b111110110010: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h8; 
end

 10'b111110110011: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h1; 
fourth_addr =4'h9; 
end

 10'b111110110100: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h0; 
end

 10'b111110110101: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h1; 
end

 10'b111110110110: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h2; 
end

 10'b111110110111: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h3; 
end

 10'b111110111000: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h4; 
end

 10'b111110111001: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h5; 
end

 10'b111110111010: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h6; 
end

 10'b111110111011: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h7; 
end

 10'b111110111100: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h8; 
end

 10'b111110111101: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h2; 
fourth_addr =4'h9; 
end

 10'b111110111110: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h0; 
end

 10'b111110111111: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h1; 
end

 10'b111111000000: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h2; 
end

 10'b111111000001: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h3; 
end

 10'b111111000010: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h4; 
end

 10'b111111000011: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h5; 
end

 10'b111111000100: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h6; 
end

 10'b111111000101: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h7; 
end

 10'b111111000110: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h8; 
end

 10'b111111000111: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h3; 
fourth_addr =4'h9; 
end

 10'b111111001000: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h0; 
end

 10'b111111001001: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h1; 
end

 10'b111111001010: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h2; 
end

 10'b111111001011: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h3; 
end

 10'b111111001100: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h4; 
end

 10'b111111001101: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h5; 
end

 10'b111111001110: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h6; 
end

 10'b111111001111: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h7; 
end

 10'b111111010000: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h8; 
end

 10'b111111010001: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h4; 
fourth_addr =4'h9; 
end

 10'b111111010010: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h0; 
end

 10'b111111010011: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h1; 
end

 10'b111111010100: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h2; 
end

 10'b111111010101: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h3; 
end

 10'b111111010110: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h4; 
end

 10'b111111010111: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h5; 
end

 10'b111111011000: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h6; 
end

 10'b111111011001: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h7; 
end

 10'b111111011010: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h8; 
end

 10'b111111011011: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h5; 
fourth_addr =4'h9; 
end

 10'b111111011100: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h0; 
end

 10'b111111011101: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h1; 
end

 10'b111111011110: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h2; 
end

 10'b111111011111: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h3; 
end

 10'b111111100000: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h4; 
end

 10'b111111100001: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h5; 
end

 10'b111111100010: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h6; 
end

 10'b111111100011: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h7; 
end

 10'b111111100100: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h8; 
end

 10'b111111100101: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h6; 
fourth_addr =4'h9; 
end

 10'b111111100110: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h0; 
end

 10'b111111100111: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h1; 
end

 10'b111111101000: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h2; 
end

 10'b111111101001: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h3; 
end

 10'b111111101010: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h4; 
end

 10'b111111101011: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h5; 
end

 10'b111111101100: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h6; 
end

 10'b111111101101: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h7; 
end

 10'b111111101110: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h8; 
end

 10'b111111101111: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h7; 
fourth_addr =4'h9; 
end

 10'b111111110000: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h0; 
end

 10'b111111110001: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h1; 
end

 10'b111111110010: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h2; 
end

 10'b111111110011: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h3; 
end

 10'b111111110100: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h4; 
end

 10'b111111110101: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h5; 
end

 10'b111111110110: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h6; 
end

 10'b111111110111: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h7; 
end

 10'b111111111000: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h8; 
end

 10'b111111111001: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h8; 
fourth_addr =4'h9; 
end

 10'b111111111010: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h0; 
end

 10'b111111111011: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h1; 
end

 10'b111111111100: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h2; 
end

 10'b111111111101: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h3; 
end

 10'b111111111110: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h4; 
end

 10'b111111111111: begin
first_addr = 4'h4; 
second_addr = 4'h0; 
third_addr = 4'h9; 
fourth_addr =4'h5; 
end
endcase
end
endmodule