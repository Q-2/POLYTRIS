
module labfinalsoc (
	clk_clk,
	generation_export_export,
	hex_digits_export,
	key_external_connection_export,
	keyboard_input_new_signal,
	keycode_export,
	leds_export,
	reset_reset_n,
	sdram_clk_clk,
	sdram_wire_addr,
	sdram_wire_ba,
	sdram_wire_cas_n,
	sdram_wire_cke,
	sdram_wire_cs_n,
	sdram_wire_dq,
	sdram_wire_dqm,
	sdram_wire_ras_n,
	sdram_wire_we_n,
	spi0_MISO,
	spi0_MOSI,
	spi0_SCLK,
	spi0_SS_n,
	usb_gpx_export,
	usb_irq_export,
	usb_rst_export,
	vga_port_blue,
	vga_port_green,
	vga_port_red,
	vga_port_hs,
	vga_port_vs,
	generator_flag_new_signal,
	game_piece_new_signal,
	random_noise_new_signal,
	piece_export_export,
	noise_export_export);	

	input		clk_clk;
	input	[7:0]	generation_export_export;
	output	[15:0]	hex_digits_export;
	input	[1:0]	key_external_connection_export;
	input	[7:0]	keyboard_input_new_signal;
	output	[7:0]	keycode_export;
	output	[13:0]	leds_export;
	input		reset_reset_n;
	output		sdram_clk_clk;
	output	[12:0]	sdram_wire_addr;
	output	[1:0]	sdram_wire_ba;
	output		sdram_wire_cas_n;
	output		sdram_wire_cke;
	output		sdram_wire_cs_n;
	inout	[15:0]	sdram_wire_dq;
	output	[1:0]	sdram_wire_dqm;
	output		sdram_wire_ras_n;
	output		sdram_wire_we_n;
	input		spi0_MISO;
	output		spi0_MOSI;
	output		spi0_SCLK;
	output		spi0_SS_n;
	input		usb_gpx_export;
	input		usb_irq_export;
	output		usb_rst_export;
	output	[3:0]	vga_port_blue;
	output	[3:0]	vga_port_green;
	output	[3:0]	vga_port_red;
	output		vga_port_hs;
	output		vga_port_vs;
	output	[7:0]	generator_flag_new_signal;
	input	[15:0]	game_piece_new_signal;
	input	[15:0]	random_noise_new_signal;
	output	[15:0]	piece_export_export;
	output	[15:0]	noise_export_export;
endmodule
