module font_rom ( input [7:0]	addr,
		  output [15:0]	data
		);

	parameter ADDR_WIDTH = 8;
   parameter DATA_WIDTH =  16;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-11][DATA_WIDTH-1:0] ROM = {
        // code x00
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b0000000000000000, // 04
        16'b0000000000000000, // 05
        16'b0000000000000000, // 06
        16'b0000000000000000, // 07
        16'b0000000000000000, // 08
        16'b0000000000000000, // 09
        16'b0000000000000000, // 0a
        16'b0000000000000000, // 0b
        16'b0000000000000000, // 0c
        16'b0000000000000000, // 0d
        16'b0000000000000000, // 0e
        16'b0000000000000000, // 0f
        // code x01
        16'b0000000000000000, // 10
        16'b0000000000000000, // 11
        16'b0000000000000000, // 12
        16'b0000000000000000, // 13
        16'b0000000000000000, // 14
        16'b0000000000000000, // 15
        16'b0000000000000000, // 16
        16'b0000000000000000, // 17
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
        // code x02
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b0011111111110000, // 04 *****
        16'b0011111111110000, // 05
        16'b1111000000111100, // 06 **   **
        16'b1111000000111100, // 07
        16'b1111000000111100, // 08 **   **
        16'b1111000000111100, // 09
        16'b1111000011111100, // 0a **  ***
        16'b1111000011111100, // 0b
        16'b1111001111111100, // 0c ** ****
        16'b1111001111111100, // 0d
        16'b1111111100111100, // 0e **** **
        16'b1111111100111100, // 0f
        // code x03
        16'b1111110000111100, // 10 ***  **
        16'b1111110000111100, // 11
        16'b1111000000111100, // 12 **   **
        16'b1111000000111100, // 13
        16'b1111000000111100, // 14 **   **
        16'b1111000000111100, // 15
        16'b0011111111110000, // 16  *****
        16'b0011111111110000, // 17
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x04
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b0000001111000000, // 04
        16'b0000001111000000, // 05
        16'b0000111111000000, // 06
        16'b0000111111000000, // 07
        16'b0011111111000000, // 08    **
        16'b0011111111000000, // 09
        16'b0000001111000000, // 0a   ***
        16'b0000001111000000, // 0b
        16'b0000001111000000, // 0c  ****
        16'b0000001111000000, // 0d
        16'b0000001111000000, // 0e    **
        16'b0000001111000000, // 0f
         // code x05
        16'b0000001111000000, // 10   **
        16'b0000001111000000, // 11
        16'b0000001111000000, // 12   **
        16'b0000001111000000, // 13
        16'b0000001111000000, // 14    **
        16'b0000001111000000, // 15
        16'b0011111111111100, // 16   **
        16'b0011111111111100, // 17
        16'b0000000000000000, // 18   **
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a ******
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x06
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b0011111111110000, // 04 *****
        16'b0011111111110000, // 05
        16'b1111000000111100, // 06 **   **
        16'b1111000000111100, // 07
        16'b0000000000111100, // 08      **
        16'b0000000000111100, // 09
        16'b0000000011110000, // 0a     **
        16'b0000000011110000, // 0b
        16'b0000001111000000, // 0c    **
        16'b0000001111000000, // 0d
        16'b0000111100000000, // 0e   **
        16'b0000111100000000, // 0f
         // code x07
        16'b0011110000000000, // 10 **
        16'b0011110000000000, // 11
        16'b1111000000000000, // 12**
        16'b1111000000000000, // 13
        16'b1111000000111100, // 14 **   **
        16'b1111000000111100, // 15
        16'b1111111111111100, // 16*******
        16'b1111111111111100, // 17
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x08
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b0011111111110000, // 04 *****
        16'b0011111111110000, // 05
        16'b1111000000111100, // 06 **   **
        16'b1111000000111100, // 07
        16'b0000000000111100, // 08      **
        16'b0000000000111100, // 09
        16'b0000000000111100, // 0a      **
        16'b0000000000111100, // 0b
        16'b0000111111110000, // 0c   ****
        16'b0000111111110000, // 0d
        16'b0000000000111100, // 0e      **
        16'b0000000000111100, // 0f
         // code x09
        16'b0000000000111100, // 10     **
        16'b0000000000111100, // 11
        16'b0000000000111100, // 12     **
        16'b0000000000111100, // 13
        16'b1111000000111100, // 14 **   **
        16'b1111000000111100, // 15
        16'b0011111111110000, // 16 *****
        16'b0011111111110000, // 17
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x0a
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b0000000011110000, // 04    **
        16'b0000000011110000, // 05
        16'b0000001111110000, // 06    ***
        16'b0000001111110000, // 07
        16'b0000111111110000, // 08   ****
        16'b0000111111110000, // 09
        16'b0011110011110000, // 0a  ** **
        16'b0011110011110000, // 0b
        16'b1111000011110000, // 0c **  **
        16'b1111000011110000, // 0d
        16'b1111111111111100, // 0e *******
        16'b1111111111111100, // 0f
         // code x0b
        16'b0000000011110000, // 10    **
        16'b0000000011110000, // 11
        16'b0000000011110000, // 12    **
        16'b0000000011110000, // 13
        16'b0000000011110000, // 14     **
        16'b0000000011110000, // 15
        16'b0000001111111100, // 16   ****
        16'b0000001111111100, // 17
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x0c
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b1111111111111100, // 04
        16'b1111111111111100, // 05
        16'b1111000000000000, // 06
        16'b1111000000000000, // 07
        16'b1111000000000000, // 08
        16'b1111000000000000, // 09
        16'b1111000000000000, // 0a
        16'b1111000000000000, // 0b
        16'b1111111111110000, // 0c
        16'b1111111111110000, // 0d
        16'b0000000000111100, // 0e
        16'b0000000000111100, // 0f
         // code x0d
        16'b0000000000111100, // 10
        16'b0000000000111100, // 11
        16'b0000000000111100, // 12
        16'b0000000000111100, // 13
        16'b1111000000111100, // 14
        16'b1111000000111100, // 15
        16'b0011111111110000, // 16
        16'b0011111111110000, // 17
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x0e
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b0000111111000000, // 04  ***
        16'b0000111111000000, // 05  ***
        16'b0011110000000000, // 06 **
        16'b0011110000000000, // 07 **
        16'b1111000000000000, // 08 **
        16'b1111000000000000, // 09 **
        16'b1111000000000000, // 0a **
        16'b1111000000000000, // 0b **
        16'b1111111111110000, // 0c ******
        16'b1111111111110000, // 0d ******
        16'b1111000000111100, // 0e **   **
        16'b1111000000111100, // 0f **   **
         // code x0f
        16'b1111000000111100, // 10 **   **
        16'b1111000000111100, // 11 **   **
        16'b1111000000111100, // 12 **   **
        16'b1111000000111100, // 13 **   **
        16'b1111000000111100, // 14 **   **
        16'b1111000000111100, // 15 **   **
        16'b0011111111110000, // 16  *****
        16'b0011111111110000, // 17  *****
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x10
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b1111111111111100, // 04*******
        16'b1111111111111100, // 05*******
        16'b1111000000111100, // 06**   **
        16'b1111000000111100, // 07**   **
        16'b0000000000111100, // 08      **
        16'b0000000000111100, // 09      **
        16'b0000000000111100, // 0a      **
        16'b0000000000111100, // 0b      **
        16'b0000000011110000, // 0c     **
        16'b0000000011110000, // 0d     **
        16'b0000001111000000, // 0e    **
        16'b0000001111000000, // 0f    **
         // code x11
        16'b0000111100000000, // 10   **
        16'b0000111100000000, // 11   **
        16'b0000111100000000, // 12   **
        16'b0000111100000000, // 13   **
        16'b0000111100000000, // 14   **
        16'b0000111100000000, // 15   **
        16'b0000111100000000, // 16   **
        16'b0000111100000000, // 17   **
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x12
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b0011111111110000, // 04 *****
        16'b0011111111110000, // 05 *****
        16'b1111000000111100, // 06**   **
        16'b1111000000111100, // 07**   **
        16'b1111000000111100, // 08 **   **
        16'b1111000000111100, // 09 **   **
        16'b1111000000111100, // 0a **   **
        16'b1111000000111100, // 0b **   **
        16'b0011111111110000, // 0c  *****
        16'b0011111111110000, // 0d  *****
        16'b1111000000111100, // 0e **   **
        16'b1111000000111100, // 0f **   **
         // code x13
        16'b1111000000111100, // 10 **   **
        16'b1111000000111100, // 11 **   **
        16'b1111000000111100, // 12 **   **
        16'b1111000000111100, // 13 **   **
        16'b1111000000111100, // 14 **   **
        16'b1111000000111100, // 15 **   **
        16'b0011111111110000, // 16  *****
        16'b0011111111110000, // 17  *****
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x14
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b0011111111110000, // 04 *****
        16'b0011111111110000, // 05 *****
        16'b1111000000111100, // 06**   **
        16'b1111000000111100, // 07**   **
        16'b1111000000111100, // 08 **   **
        16'b1111000000111100, // 09 **   **
        16'b1111000000111100, // 0a **   **
        16'b1111000000111100, // 0b **   **
        16'b0011111111111100, // 0c  ******
        16'b0011111111111100, // 0d  ******
        16'b0000000000111100, // 0e      **
        16'b0000000000111100, // 0f      **
         // code x15
        16'b0000000000111100, // 10      **
        16'b0000000000111100, // 11      **
        16'b0000000000111100, // 12      **
        16'b0000000000111100, // 13      **
        16'b0000000011110000, // 14     **
        16'b0000000011110000, // 15     **
        16'b0011111111000000, // 16  ****
        16'b0011111111000000, // 17  ****
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x16
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b0000001100000000, // 04   *
        16'b0000001100000000, // 05   *
        16'b0000111111000000, // 06  ***
        16'b0000111111000000, // 07  ***
        16'b0011110011110000, // 08  ** **
        16'b0011110011110000, // 09  ** **
        16'b1111000000111100, // 0a **   **
        16'b1111000000111100, // 0b **   **
        16'b1111000000111100, // 0c **   **
        16'b1111000000111100, // 0d **   **
        16'b1111111111111100, // 0e *******
        16'b1111111111111100, // 0f *******
         // code x17
        16'b1111000000111100, // 10 **   **
        16'b1111000000111100, // 11 **   **
        16'b1111000000111100, // 12 **   **
        16'b1111000000111100, // 13 **   **
        16'b1111000000111100, // 14 **   **
        16'b1111000000111100, // 15 **   **
        16'b1111000000111100, // 16 **   **
        16'b1111000000111100, // 17 **   **
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x18
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b0000111111110000, // 04  ****
        16'b0000111111110000, // 05  ****
        16'b0011110000111100, // 06 **  **
        16'b0011110000111100, // 07 **  **
        16'b1111000000001100, // 08 **    *
        16'b1111000000001100, // 09 **    *
        16'b1111000000000000, // 0a **
        16'b1111000000000000, // 0b **
        16'b1111000000000000, // 0c **
        16'b1111000000000000, // 0d **
        16'b1111000000000000, // 0e **
        16'b1111000000000000, // 0f **
         // code x19
        16'b1111000000000000, // 10 **
        16'b1111000000000000, // 11 **
        16'b1111000000001100, // 12 **    *
        16'b1111000000001100, // 13 **    *
        16'b0011110000111100, // 14  **  **
        16'b0011110000111100, // 15  **  **
        16'b0000111111110000, // 16   ****
        16'b0000111111110000, // 17   ****
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x1a
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b1111111111111100, // 04*******
        16'b1111111111111100, // 05*******
        16'b0011110000111100, // 06 **  **
        16'b0011110000111100, // 07 **  **
        16'b0011110000001100, // 08  **   *
        16'b0011110000001100, // 09  **   *
        16'b0011110011000000, // 0a  ** *
        16'b0011110011000000, // 0b  ** *
        16'b0011111111000000, // 0c  ****
        16'b0011111111000000, // 0d  ****
        16'b0011110011000000, // 0e  ** *
        16'b0011110011000000, // 0f  ** *
         // code x1b
        16'b0011110000000000, // 10  **
        16'b0011110000000000, // 11  **
        16'b0011110000001100, // 12  **   *
        16'b0011110000001100, // 13  **   *
        16'b0011110000111100, // 14  **  **
        16'b0011110000111100, // 15  **  **
        16'b1111111111111100, // 16 *******
        16'b1111111111111100, // 17 *******
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x1c
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b0000111111110000, // 04  ****
        16'b0000111111110000, // 05  ****
        16'b0000001111000000, // 06   **
        16'b0000001111000000, // 07   **
        16'b0000001111000000, // 08    **
        16'b0000001111000000, // 09    **
        16'b0000001111000000, // 0a    **
        16'b0000001111000000, // 0b    **
        16'b0000001111000000, // 0c    **
        16'b0000001111000000, // 0d    **
        16'b0000001111000000, // 0e    **
        16'b0000001111000000, // 0f    **
         // code x1d
        16'b0000001111000000, // 10    **
        16'b0000001111000000, // 11    **
        16'b0000001111000000, // 12    **
        16'b0000001111000000, // 13    **
        16'b0000001111000000, // 14    **
        16'b0000001111000000, // 15    **
        16'b0000111111110000, // 16   ****
        16'b0000111111110000, // 17   ****
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x1e
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b1111111100000000, // 04****
        16'b1111111100000000, // 05****
        16'b0011110000000000, // 06 **
        16'b0011110000000000, // 07 **
        16'b0011110000000000, // 08  **
        16'b0011110000000000, // 09  **
        16'b0011110000000000, // 0a  **
        16'b0011110000000000, // 0b  **
        16'b0011110000000000, // 0c  **
        16'b0011110000000000, // 0d  **
        16'b0011110000000000, // 0e  **
        16'b0011110000000000, // 0f  **
         // code x1f
        16'b0011110000000000, // 10  **
        16'b0011110000000000, // 11  **
        16'b0011110000001100, // 12  **   *
        16'b0011110000001100, // 13  **   *
        16'b0011110000111100, // 14  **  **
        16'b0011110000111100, // 15  **  **
        16'b1111111111111100, // 16 *******
        16'b1111111111111100, // 17 *******
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x20
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b1111000000111100, // 04**   **
        16'b1111000000111100, // 05**   **
        16'b1111110000111100, // 06***  **
        16'b1111110000111100, // 07***  **
        16'b1111111100111100, // 08 **** **
        16'b1111111100111100, // 09 **** **
        16'b1111111111111100, // 0a *******
        16'b1111111111111100, // 0b *******
        16'b1111001111111100, // 0c ** ****
        16'b1111001111111100, // 0d ** ****
        16'b1111000011111100, // 0e **  ***
        16'b1111000011111100, // 0f **  ***
         // code x21
        16'b1111000000111100, // 10 **   **
        16'b1111000000111100, // 11 **   **
        16'b1111000000111100, // 12 **   **
        16'b1111000000111100, // 13 **   **
        16'b1111000000111100, // 14 **   **
        16'b1111000000111100, // 15 **   **
        16'b1111000000111100, // 16 **   **
        16'b1111000000111100, // 17 **   **
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x22
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b0011111111110000, // 04 *****
        16'b0011111111110000, // 05 *****
        16'b1111000000111100, // 06**   **
        16'b1111000000111100, // 07**   **
        16'b1111000000111100, // 08 **   **
        16'b1111000000111100, // 09 **   **
        16'b1111000000111100, // 0a **   **
        16'b1111000000111100, // 0b **   **
        16'b1111000000111100, // 0c **   **
        16'b1111000000111100, // 0d **   **
        16'b1111000000111100, // 0e **   **
        16'b1111000000111100, // 0f **   **
         // code x23
        16'b1111000000111100, // 10 **   **
        16'b1111000000111100, // 11 **   **
        16'b1111000000111100, // 12 **   **
        16'b1111000000111100, // 13 **   **
        16'b1111000000111100, // 14 **   **
        16'b1111000000111100, // 15 **   **
        16'b0011111111110000, // 16  *****
        16'b0011111111110000, // 17  *****
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x24
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b1111111111110000, // 04******
        16'b1111111111110000, // 05******
        16'b0011110000111100, // 06 **  **
        16'b0011110000111100, // 07 **  **
        16'b0011110000111100, // 08  **  **
        16'b0011110000111100, // 09  **  **
        16'b0011110000111100, // 0a  **  **
        16'b0011110000111100, // 0b  **  **
        16'b0011111111110000, // 0c  *****
        16'b0011111111110000, // 0d  *****
        16'b0011110011110000, // 0e  ** **
        16'b0011110011110000, // 0f  ** **
         // code x25
        16'b0011110000111100, // 10  **  **
        16'b0011110000111100, // 11  **  **
        16'b0011110000111100, // 12  **  **
        16'b0011110000111100, // 13  **  **
        16'b0011110000111100, // 14  **  **
        16'b0011110000111100, // 15  **  **
        16'b1111110000111100, // 16 ***  **
        16'b1111110000111100, // 17 ***  **
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x26
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b0011111111110000, // 04 *****
        16'b0011111111110000, // 05 *****
        16'b1111000000111100, // 06**   **
        16'b1111000000111100, // 07**   **
        16'b1111000000111100, // 08 **   **
        16'b1111000000111100, // 09 **   **
        16'b0011110000000000, // 0a  **
        16'b0011110000000000, // 0b  **
        16'b0000111111000000, // 0c   ***
        16'b0000111111000000, // 0d   ***
        16'b0000000011110000, // 0e     **
        16'b0000000011110000, // 0f     **
         // code x27
        16'b0000000000111100, // 10      **
        16'b0000000000111100, // 11      **
        16'b1111000000111100, // 12 **   **
        16'b1111000000111100, // 13 **   **
        16'b1111000000111100, // 14 **   **
        16'b1111000000111100, // 15 **   **
        16'b0011111111110000, // 16  *****
        16'b0011111111110000, // 17  *****
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x28
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b1111111111111111, // 04********
        16'b1111111111111111, // 05********
        16'b1111001111001111, // 06** ** **
        16'b1111001111001111, // 07** ** **
        16'b1100001111000011, // 08 *  **  *
        16'b1100001111000011, // 09 *  **  *
        16'b0000001111000000, // 0a    **
        16'b0000001111000000, // 0b    **
        16'b0000001111000000, // 0c    **
        16'b0000001111000000, // 0d    **
        16'b0000001111000000, // 0e    **
        16'b0000001111000000, // 0f    **
         // code x29
        16'b0000001111000000, // 10    **
        16'b0000001111000000, // 11    **
        16'b0000001111000000, // 12    **
        16'b0000001111000000, // 13    **
        16'b0000001111000000, // 14    **
        16'b0000001111000000, // 15    **
        16'b0000111111110000, // 16   ****
        16'b0000111111110000, // 17   ****
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x2a
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b1111000000001111, // 04**    **
        16'b1111000000001111, // 05**    **
        16'b1111000000001111, // 06**    **
        16'b1111000000001111, // 07**    **
        16'b1111000000001111, // 08 **    **
        16'b1111000000001111, // 09 **    **
        16'b1111000000001111, // 0a **    **
        16'b1111000000001111, // 0b **    **
        16'b1111000000001111, // 0c **    **
        16'b1111000000001111, // 0d **    **
        16'b1111000000001111, // 0e **    **
        16'b1111000000001111, // 0f **    **
         // code x2b
        16'b1111000000001111, // 10 **    **
        16'b1111000000001111, // 11 **    **
        16'b0011110000111100, // 12  **  **
        16'b0011110000111100, // 13  **  **
        16'b0000111111110000, // 14   ****
        16'b0000111111110000, // 15   ****
        16'b0000001111000000, // 16    **
        16'b0000001111000000, // 17    **
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f
         // code x2c
        16'b0000000000000000, // 00
        16'b0000000000000000, // 01
        16'b0000000000000000, // 02
        16'b0000000000000000, // 03
        16'b1111000000001111, // 04**    **
        16'b1111000000001111, // 05**    **
        16'b1111000000001111, // 06**    **
        16'b1111000000001111, // 07**    **
        16'b0011110000111100, // 08  **  **
        16'b0011110000111100, // 09  **  **
        16'b0000111111110000, // 0a   ****
        16'b0000111111110000, // 0b   ****
        16'b0000001111000000, // 0c    **
        16'b0000001111000000, // 0d    **
        16'b0000001111000000, // 0e    **
        16'b0000001111000000, // 0f    **
         // code x2d
        16'b0000111111110000, // 10   ****
        16'b0000111111110000, // 11   ****
        16'b0011110000111100, // 12  **  **
        16'b0011110000111100, // 13  **  **
        16'b1111000000001111, // 14 **    **
        16'b1111000000001111, // 15 **    **
        16'b1111000000001111, // 16 **    **
        16'b1111000000001111, // 17 **    **
        16'b0000000000000000, // 18
        16'b0000000000000000, // 19
        16'b0000000000000000, // 1a
        16'b0000000000000000, // 1b
        16'b0000000000000000, // 1c
        16'b0000000000000000, // 1d
        16'b0000000000000000, // 1e
        16'b0000000000000000, // 1f

        };

	assign data = ROM[addr];

endmodule  