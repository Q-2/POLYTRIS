module drawing(
    input [5:0] SPRITE_ADDR,
	output [31:0] SPRITE_DATA
    );

    parameter ADDR_WIDTH = 6;
    parameter DATA_WIDTH =  32;
//	logic [ADDR_WIDTH-1:0] addr_reg;    //never used
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
        // blank block      x00
        32'b10101010101010101010101010101010, // 0
        32'b10101010101010101010101010101010, // 1
        32'b10101010101010101010101010101010, // 2
        32'b10101010101010101010101010101010, // 3
        32'b10101010101010101010101010101010, // 4
        32'b10101010101010101010101010101010, // 5
        32'b10101010101010101010101010101010, // 6
        32'b10101010101010101010101010101010, // 7
        32'b10101010101010101010101010101010, // 8
        32'b10101010101010101010101010101010, // 9
        32'b10101010101010101010101010101010, // a
        32'b10101010101010101010101010101010, // b
        32'b10101010101010101010101010101010, // c
        32'b10101010101010101010101010101010, // d
        32'b10101010101010101010101010101010, // e
        32'b10101010101010101010101010101010, // f
        // block style 1    x01
        32'b00000000000000000000000000000000, // 0
        32'b00000000000000000000000000000000, // 1
        32'b00001111111100000000000000000000, // 2
        32'b00001111111100000000000000000000, // 3
        32'b00001111000000000000000000000000, // 4
        32'b00001111000000000000000000000000, // 5
        32'b00000000000000000000000000000000, // 6
        32'b00000000000000000000000000000000, // 7
        32'b00000000000000000000000000000000, // 8
        32'b00000000000000000000000000000000, // 9
        32'b00000000000000000000000000000000, // a
        32'b00000000000000000000000000000000, // b
        32'b00000000000000000000000000000000, // c
        32'b00000000000000000000000000000000, // d
        32'b00000000000000000000000000000000, // e
        32'b00000000000000000000000000000000, // f
         // block style 2   x02
        32'b01010101010101010101010101010101, // 0
        32'b01010101010101010101010101010101, // 1
        32'b01011111111101010101010101010101, // 2
        32'b01011111111101010101010101010101, // 3
        32'b01011111010101010101010101010101, // 4
        32'b01011111010101010101010101010101, // 5
        32'b01010101010101010101010101010101, // 6
        32'b01010101010101010101010101010101, // 7
        32'b01010101010101010101010101010101, // 8
        32'b01010101010101010101010101010101, // 9
        32'b01010101010101010101010101010101, // a
        32'b01010101010101010101010101010101, // b
        32'b01010101010101010101010101010101, // c
        32'b01010101010101010101010101010101, // d
        32'b01010101010101010101010101010101, // e
        32'b01010101010101010101010101010101, // f
         // block style 3   x03
        32'b00000000000000000000000000000000, // 0
        32'b00000000000000000000000000000000, // 1
        32'b00001111111111111111111111110000, // 2
        32'b00001111111111111111111111110000, // 3
        32'b00001111111111111111111111110000, // 4
        32'b00001111111111111111111111110000, // 5
        32'b00001111111111111111111111110000, // 6
        32'b00001111111111111111111111110000, // 7
        32'b00001111111111111111111111110000, // 8
        32'b00001111111111111111111111110000, // 9
        32'b00001111111111111111111111110000, // a
        32'b00001111111111111111111111110000, // b
        32'b00001111111111111111111111110000, // c
        32'b00001111111111111111111111110000, // d
        32'b00000000000000000000000000000000, // e
        32'b00000000000000000000000000000000, // f

        };

	assign SPRITE_DATA = ROM[SPRITE_ADDR]; 

endmodule
