// labfinalsoc.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module labfinalsoc (
		input  wire        clk_clk,                        //                     clk.clk
		input  wire [15:0] game_piece_new_signal,          //              game_piece.new_signal
		input  wire [7:0]  generation_export_export,       //       generation_export.export
		output wire [7:0]  generator_flag_new_signal,      //          generator_flag.new_signal
		output wire [15:0] hex_digits_export,              //              hex_digits.export
		input  wire [1:0]  key_external_connection_export, // key_external_connection.export
		input  wire [7:0]  keyboard_input_new_signal,      //          keyboard_input.new_signal
		output wire [7:0]  keycode_export,                 //                 keycode.export
		output wire [13:0] leds_export,                    //                    leds.export
		output wire [15:0] noise_export_export,            //            noise_export.export
		output wire [15:0] piece_export_export,            //            piece_export.export
		input  wire [15:0] random_noise_new_signal,        //            random_noise.new_signal
		input  wire        reset_reset_n,                  //                   reset.reset_n
		output wire        sdram_clk_clk,                  //               sdram_clk.clk
		output wire [12:0] sdram_wire_addr,                //              sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                  //                        .ba
		output wire        sdram_wire_cas_n,               //                        .cas_n
		output wire        sdram_wire_cke,                 //                        .cke
		output wire        sdram_wire_cs_n,                //                        .cs_n
		inout  wire [15:0] sdram_wire_dq,                  //                        .dq
		output wire [1:0]  sdram_wire_dqm,                 //                        .dqm
		output wire        sdram_wire_ras_n,               //                        .ras_n
		output wire        sdram_wire_we_n,                //                        .we_n
		input  wire        spi0_MISO,                      //                    spi0.MISO
		output wire        spi0_MOSI,                      //                        .MOSI
		output wire        spi0_SCLK,                      //                        .SCLK
		output wire        spi0_SS_n,                      //                        .SS_n
		input  wire        usb_gpx_export,                 //                 usb_gpx.export
		input  wire        usb_irq_export,                 //                 usb_irq.export
		output wire        usb_rst_export,                 //                 usb_rst.export
		output wire [3:0]  vga_port_blue,                  //                vga_port.blue
		output wire [3:0]  vga_port_green,                 //                        .green
		output wire [3:0]  vga_port_red,                   //                        .red
		output wire        vga_port_hs,                    //                        .hs
		output wire        vga_port_vs                     //                        .vs
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                                       // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                                    // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                                    // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [27:0] nios2_gen2_0_data_master_address;                                        // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                                     // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                           // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                                          // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                                      // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                                // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                             // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [27:0] nios2_gen2_0_instruction_master_address;                                 // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                                    // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                  // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;               // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                 // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_chipselect; // mm_interconnect_0:VGA_text_mode_controller_0_avalon_mm_slave_chipselect -> VGA_text_mode_controller_0:AVL_CS
	wire  [31:0] mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_readdata;   // VGA_text_mode_controller_0:AVL_READDATA -> mm_interconnect_0:VGA_text_mode_controller_0_avalon_mm_slave_readdata
	wire  [11:0] mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_address;    // mm_interconnect_0:VGA_text_mode_controller_0_avalon_mm_slave_address -> VGA_text_mode_controller_0:AVL_ADDR
	wire         mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_read;       // mm_interconnect_0:VGA_text_mode_controller_0_avalon_mm_slave_read -> VGA_text_mode_controller_0:AVL_READ
	wire   [3:0] mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_byteenable; // mm_interconnect_0:VGA_text_mode_controller_0_avalon_mm_slave_byteenable -> VGA_text_mode_controller_0:AVL_BYTE_EN
	wire         mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_write;      // mm_interconnect_0:VGA_text_mode_controller_0_avalon_mm_slave_write -> VGA_text_mode_controller_0:AVL_WRITE
	wire  [31:0] mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_writedata;  // mm_interconnect_0:VGA_text_mode_controller_0_avalon_mm_slave_writedata -> VGA_text_mode_controller_0:AVL_WRITEDATA
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;                   // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;                    // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;                 // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;              // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;              // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;                  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;                     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;               // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;                    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;                // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;                           // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;                            // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                               // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                              // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;                          // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                        // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                          // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [1:0] mm_interconnect_0_onchip_memory2_0_s1_address;                           // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                        // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                             // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                         // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                             // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                                   // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                     // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                  // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                      // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                         // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                   // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                        // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                    // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_keycode_s1_chipselect;                                 // mm_interconnect_0:keycode_s1_chipselect -> keycode:chipselect
	wire  [31:0] mm_interconnect_0_keycode_s1_readdata;                                   // keycode:readdata -> mm_interconnect_0:keycode_s1_readdata
	wire   [1:0] mm_interconnect_0_keycode_s1_address;                                    // mm_interconnect_0:keycode_s1_address -> keycode:address
	wire         mm_interconnect_0_keycode_s1_write;                                      // mm_interconnect_0:keycode_s1_write -> keycode:write_n
	wire  [31:0] mm_interconnect_0_keycode_s1_writedata;                                  // mm_interconnect_0:keycode_s1_writedata -> keycode:writedata
	wire  [31:0] mm_interconnect_0_usb_irq_s1_readdata;                                   // usb_irq:readdata -> mm_interconnect_0:usb_irq_s1_readdata
	wire   [1:0] mm_interconnect_0_usb_irq_s1_address;                                    // mm_interconnect_0:usb_irq_s1_address -> usb_irq:address
	wire  [31:0] mm_interconnect_0_usb_gpx_s1_readdata;                                   // usb_gpx:readdata -> mm_interconnect_0:usb_gpx_s1_readdata
	wire   [1:0] mm_interconnect_0_usb_gpx_s1_address;                                    // mm_interconnect_0:usb_gpx_s1_address -> usb_gpx:address
	wire         mm_interconnect_0_hex_digits_s1_chipselect;                              // mm_interconnect_0:hex_digits_s1_chipselect -> hex_digits:chipselect
	wire  [31:0] mm_interconnect_0_hex_digits_s1_readdata;                                // hex_digits:readdata -> mm_interconnect_0:hex_digits_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_digits_s1_address;                                 // mm_interconnect_0:hex_digits_s1_address -> hex_digits:address
	wire         mm_interconnect_0_hex_digits_s1_write;                                   // mm_interconnect_0:hex_digits_s1_write -> hex_digits:write_n
	wire  [31:0] mm_interconnect_0_hex_digits_s1_writedata;                               // mm_interconnect_0:hex_digits_s1_writedata -> hex_digits:writedata
	wire         mm_interconnect_0_leds_pio_s1_chipselect;                                // mm_interconnect_0:leds_pio_s1_chipselect -> leds_pio:chipselect
	wire  [31:0] mm_interconnect_0_leds_pio_s1_readdata;                                  // leds_pio:readdata -> mm_interconnect_0:leds_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_pio_s1_address;                                   // mm_interconnect_0:leds_pio_s1_address -> leds_pio:address
	wire         mm_interconnect_0_leds_pio_s1_write;                                     // mm_interconnect_0:leds_pio_s1_write -> leds_pio:write_n
	wire  [31:0] mm_interconnect_0_leds_pio_s1_writedata;                                 // mm_interconnect_0:leds_pio_s1_writedata -> leds_pio:writedata
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                                       // key:readdata -> mm_interconnect_0:key_s1_readdata
	wire   [1:0] mm_interconnect_0_key_s1_address;                                        // mm_interconnect_0:key_s1_address -> key:address
	wire         mm_interconnect_0_timer_s1_chipselect;                                   // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                                     // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [3:0] mm_interconnect_0_timer_s1_address;                                      // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                                        // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                                    // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_usb_rst_s1_chipselect;                                 // mm_interconnect_0:usb_rst_s1_chipselect -> usb_rst:chipselect
	wire  [31:0] mm_interconnect_0_usb_rst_s1_readdata;                                   // usb_rst:readdata -> mm_interconnect_0:usb_rst_s1_readdata
	wire   [1:0] mm_interconnect_0_usb_rst_s1_address;                                    // mm_interconnect_0:usb_rst_s1_address -> usb_rst:address
	wire         mm_interconnect_0_usb_rst_s1_write;                                      // mm_interconnect_0:usb_rst_s1_write -> usb_rst:write_n
	wire  [31:0] mm_interconnect_0_usb_rst_s1_writedata;                                  // mm_interconnect_0:usb_rst_s1_writedata -> usb_rst:writedata
	wire  [31:0] mm_interconnect_0_generator_pio_s1_readdata;                             // generator_pio:readdata -> mm_interconnect_0:generator_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_generator_pio_s1_address;                              // mm_interconnect_0:generator_pio_s1_address -> generator_pio:address
	wire         mm_interconnect_0_piece_pio_s1_chipselect;                               // mm_interconnect_0:piece_pio_s1_chipselect -> piece_pio:chipselect
	wire  [31:0] mm_interconnect_0_piece_pio_s1_readdata;                                 // piece_pio:readdata -> mm_interconnect_0:piece_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_piece_pio_s1_address;                                  // mm_interconnect_0:piece_pio_s1_address -> piece_pio:address
	wire         mm_interconnect_0_piece_pio_s1_write;                                    // mm_interconnect_0:piece_pio_s1_write -> piece_pio:write_n
	wire  [31:0] mm_interconnect_0_piece_pio_s1_writedata;                                // mm_interconnect_0:piece_pio_s1_writedata -> piece_pio:writedata
	wire         mm_interconnect_0_noise_pio_s1_chipselect;                               // mm_interconnect_0:noise_pio_s1_chipselect -> noise_pio:chipselect
	wire  [31:0] mm_interconnect_0_noise_pio_s1_readdata;                                 // noise_pio:readdata -> mm_interconnect_0:noise_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_noise_pio_s1_address;                                  // mm_interconnect_0:noise_pio_s1_address -> noise_pio:address
	wire         mm_interconnect_0_noise_pio_s1_write;                                    // mm_interconnect_0:noise_pio_s1_write -> noise_pio:write_n
	wire  [31:0] mm_interconnect_0_noise_pio_s1_writedata;                                // mm_interconnect_0:noise_pio_s1_writedata -> noise_pio:writedata
	wire         mm_interconnect_0_spi_0_spi_control_port_chipselect;                     // mm_interconnect_0:spi_0_spi_control_port_chipselect -> spi_0:spi_select
	wire  [15:0] mm_interconnect_0_spi_0_spi_control_port_readdata;                       // spi_0:data_to_cpu -> mm_interconnect_0:spi_0_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_0_spi_control_port_address;                        // mm_interconnect_0:spi_0_spi_control_port_address -> spi_0:mem_addr
	wire         mm_interconnect_0_spi_0_spi_control_port_read;                           // mm_interconnect_0:spi_0_spi_control_port_read -> spi_0:read_n
	wire         mm_interconnect_0_spi_0_spi_control_port_write;                          // mm_interconnect_0:spi_0_spi_control_port_write -> spi_0:write_n
	wire  [15:0] mm_interconnect_0_spi_0_spi_control_port_writedata;                      // mm_interconnect_0:spi_0_spi_control_port_writedata -> spi_0:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                                // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                // timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                // spi_0:irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                                    // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                                          // rst_controller:reset_out -> [VGA_text_mode_controller_0:RESET, generator_pio:reset_n, mm_interconnect_0:VGA_text_mode_controller_0_RESET_reset_bridge_in_reset_reset, noise_pio:reset_n, piece_pio:reset_n]
	wire         rst_controller_001_reset_out_reset;                                      // rst_controller_001:reset_out -> [altpll_0:reset, hex_digits:reset_n, irq_mapper:reset, jtag_uart:rst_n, key:reset_n, keycode:reset_n, leds_pio:reset_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, sdram:reset_n, spi_0:reset_n, sysid_qsys_0:reset_n, timer:reset_n, usb_gpx:reset_n, usb_irq:reset_n, usb_rst:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                                  // rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                                  // nios2_gen2_0:debug_reset_request -> rst_controller_001:reset_in1

	vga_text_avl_interface vga_text_mode_controller_0 (
		.CLK            (clk_clk),                                                                 //             CLK.clk
		.RESET          (rst_controller_reset_out_reset),                                          //           RESET.reset
		.AVL_CS         (mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_chipselect), // avalon_mm_slave.chipselect
		.AVL_BYTE_EN    (mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_byteenable), //                .byteenable
		.AVL_ADDR       (mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_address),    //                .address
		.AVL_READ       (mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_read),       //                .read
		.AVL_READDATA   (mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_readdata),   //                .readdata
		.AVL_WRITE      (mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_write),      //                .write
		.AVL_WRITEDATA  (mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_writedata),  //                .writedata
		.blue           (vga_port_blue),                                                           //        VGA_port.blue
		.green          (vga_port_green),                                                          //                .green
		.red            (vga_port_red),                                                            //                .red
		.hs             (vga_port_hs),                                                             //                .hs
		.vs             (vga_port_vs),                                                             //                .vs
		.keyboard_input (keyboard_input_new_signal),                                               //        keyboard.new_signal
		.generator_flag (generator_flag_new_signal),                                               //       generator.new_signal
		.game_piece     (game_piece_new_signal),                                                   //           piece.new_signal
		.random_noise   (random_noise_new_signal)                                                  //           noise.new_signal
	);

	labfinalsoc_altpll_0 altpll_0 (
		.clk                (clk_clk),                                        //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),             // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0                 (),                                               //                    c0.clk
		.c1                 (sdram_clk_clk),                                  //                    c1.clk
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.c2                 (),                                               //           (terminated)
		.c3                 (),                                               //           (terminated)
		.c4                 (),                                               //           (terminated)
		.areset             (1'b0),                                           //           (terminated)
		.locked             (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (3'b000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	labfinalsoc_generator_pio generator_pio (
		.clk      (clk_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_generator_pio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_generator_pio_s1_readdata), //                    .readdata
		.in_port  (generation_export_export)                     // external_connection.export
	);

	labfinalsoc_hex_digits hex_digits (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_hex_digits_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_digits_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_digits_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_digits_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_digits_s1_readdata),   //                    .readdata
		.out_port   (hex_digits_export)                           // external_connection.export
	);

	labfinalsoc_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	labfinalsoc_key key (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_key_s1_address),    //                  s1.address
		.readdata (mm_interconnect_0_key_s1_readdata),   //                    .readdata
		.in_port  (key_external_connection_export)       // external_connection.export
	);

	labfinalsoc_keycode keycode (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_keycode_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keycode_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keycode_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keycode_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keycode_s1_readdata),   //                    .readdata
		.out_port   (keycode_export)                           // external_connection.export
	);

	labfinalsoc_leds_pio leds_pio (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_pio_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                               // external_connection.export
	);

	labfinalsoc_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	labfinalsoc_hex_digits noise_pio (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_noise_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_noise_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_noise_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_noise_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_noise_pio_s1_readdata),   //                    .readdata
		.out_port   (noise_export_export)                        // external_connection.export
	);

	labfinalsoc_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	labfinalsoc_hex_digits piece_pio (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_piece_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_piece_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_piece_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_piece_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_piece_pio_s1_readdata),   //                    .readdata
		.out_port   (piece_export_export)                        // external_connection.export
	);

	labfinalsoc_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	labfinalsoc_spi_0 spi_0 (
		.clk           (clk_clk),                                             //              clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                 //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_0_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_0_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_0_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_0_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_0_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_0_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver2_irq),                            //              irq.irq
		.MISO          (spi0_MISO),                                           //         external.export
		.MOSI          (spi0_MOSI),                                           //                 .export
		.SCLK          (spi0_SCLK),                                           //                 .export
		.SS_n          (spi0_SS_n)                                            //                 .export
	);

	labfinalsoc_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	labfinalsoc_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	labfinalsoc_usb_gpx usb_gpx (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_usb_gpx_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_usb_gpx_s1_readdata), //                    .readdata
		.in_port  (usb_gpx_export)                         // external_connection.export
	);

	labfinalsoc_usb_gpx usb_irq (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_usb_irq_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_usb_irq_s1_readdata), //                    .readdata
		.in_port  (usb_irq_export)                         // external_connection.export
	);

	labfinalsoc_usb_rst usb_rst (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_usb_rst_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_usb_rst_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_usb_rst_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_usb_rst_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_usb_rst_s1_readdata),   //                    .readdata
		.out_port   (usb_rst_export)                           // external_connection.export
	);

	labfinalsoc_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                                (clk_clk),                                                                 //                                              clk_0_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset               (rst_controller_001_reset_out_reset),                                      //               nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.VGA_text_mode_controller_0_RESET_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                          // VGA_text_mode_controller_0_RESET_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                             (nios2_gen2_0_data_master_address),                                        //                               nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                         (nios2_gen2_0_data_master_waitrequest),                                    //                                                       .waitrequest
		.nios2_gen2_0_data_master_byteenable                          (nios2_gen2_0_data_master_byteenable),                                     //                                                       .byteenable
		.nios2_gen2_0_data_master_read                                (nios2_gen2_0_data_master_read),                                           //                                                       .read
		.nios2_gen2_0_data_master_readdata                            (nios2_gen2_0_data_master_readdata),                                       //                                                       .readdata
		.nios2_gen2_0_data_master_write                               (nios2_gen2_0_data_master_write),                                          //                                                       .write
		.nios2_gen2_0_data_master_writedata                           (nios2_gen2_0_data_master_writedata),                                      //                                                       .writedata
		.nios2_gen2_0_data_master_debugaccess                         (nios2_gen2_0_data_master_debugaccess),                                    //                                                       .debugaccess
		.nios2_gen2_0_instruction_master_address                      (nios2_gen2_0_instruction_master_address),                                 //                        nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                  (nios2_gen2_0_instruction_master_waitrequest),                             //                                                       .waitrequest
		.nios2_gen2_0_instruction_master_read                         (nios2_gen2_0_instruction_master_read),                                    //                                                       .read
		.nios2_gen2_0_instruction_master_readdata                     (nios2_gen2_0_instruction_master_readdata),                                //                                                       .readdata
		.altpll_0_pll_slave_address                                   (mm_interconnect_0_altpll_0_pll_slave_address),                            //                                     altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                     (mm_interconnect_0_altpll_0_pll_slave_write),                              //                                                       .write
		.altpll_0_pll_slave_read                                      (mm_interconnect_0_altpll_0_pll_slave_read),                               //                                                       .read
		.altpll_0_pll_slave_readdata                                  (mm_interconnect_0_altpll_0_pll_slave_readdata),                           //                                                       .readdata
		.altpll_0_pll_slave_writedata                                 (mm_interconnect_0_altpll_0_pll_slave_writedata),                          //                                                       .writedata
		.generator_pio_s1_address                                     (mm_interconnect_0_generator_pio_s1_address),                              //                                       generator_pio_s1.address
		.generator_pio_s1_readdata                                    (mm_interconnect_0_generator_pio_s1_readdata),                             //                                                       .readdata
		.hex_digits_s1_address                                        (mm_interconnect_0_hex_digits_s1_address),                                 //                                          hex_digits_s1.address
		.hex_digits_s1_write                                          (mm_interconnect_0_hex_digits_s1_write),                                   //                                                       .write
		.hex_digits_s1_readdata                                       (mm_interconnect_0_hex_digits_s1_readdata),                                //                                                       .readdata
		.hex_digits_s1_writedata                                      (mm_interconnect_0_hex_digits_s1_writedata),                               //                                                       .writedata
		.hex_digits_s1_chipselect                                     (mm_interconnect_0_hex_digits_s1_chipselect),                              //                                                       .chipselect
		.jtag_uart_avalon_jtag_slave_address                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                   //                            jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                     //                                                       .write
		.jtag_uart_avalon_jtag_slave_read                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                      //                                                       .read
		.jtag_uart_avalon_jtag_slave_readdata                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),                  //                                                       .readdata
		.jtag_uart_avalon_jtag_slave_writedata                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),                 //                                                       .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),               //                                                       .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),                //                                                       .chipselect
		.key_s1_address                                               (mm_interconnect_0_key_s1_address),                                        //                                                 key_s1.address
		.key_s1_readdata                                              (mm_interconnect_0_key_s1_readdata),                                       //                                                       .readdata
		.keycode_s1_address                                           (mm_interconnect_0_keycode_s1_address),                                    //                                             keycode_s1.address
		.keycode_s1_write                                             (mm_interconnect_0_keycode_s1_write),                                      //                                                       .write
		.keycode_s1_readdata                                          (mm_interconnect_0_keycode_s1_readdata),                                   //                                                       .readdata
		.keycode_s1_writedata                                         (mm_interconnect_0_keycode_s1_writedata),                                  //                                                       .writedata
		.keycode_s1_chipselect                                        (mm_interconnect_0_keycode_s1_chipselect),                                 //                                                       .chipselect
		.leds_pio_s1_address                                          (mm_interconnect_0_leds_pio_s1_address),                                   //                                            leds_pio_s1.address
		.leds_pio_s1_write                                            (mm_interconnect_0_leds_pio_s1_write),                                     //                                                       .write
		.leds_pio_s1_readdata                                         (mm_interconnect_0_leds_pio_s1_readdata),                                  //                                                       .readdata
		.leds_pio_s1_writedata                                        (mm_interconnect_0_leds_pio_s1_writedata),                                 //                                                       .writedata
		.leds_pio_s1_chipselect                                       (mm_interconnect_0_leds_pio_s1_chipselect),                                //                                                       .chipselect
		.nios2_gen2_0_debug_mem_slave_address                         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),                  //                           nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),                    //                                                       .write
		.nios2_gen2_0_debug_mem_slave_read                            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),                     //                                                       .read
		.nios2_gen2_0_debug_mem_slave_readdata                        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),                 //                                                       .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),                //                                                       .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                      (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),               //                                                       .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),              //                                                       .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),              //                                                       .debugaccess
		.noise_pio_s1_address                                         (mm_interconnect_0_noise_pio_s1_address),                                  //                                           noise_pio_s1.address
		.noise_pio_s1_write                                           (mm_interconnect_0_noise_pio_s1_write),                                    //                                                       .write
		.noise_pio_s1_readdata                                        (mm_interconnect_0_noise_pio_s1_readdata),                                 //                                                       .readdata
		.noise_pio_s1_writedata                                       (mm_interconnect_0_noise_pio_s1_writedata),                                //                                                       .writedata
		.noise_pio_s1_chipselect                                      (mm_interconnect_0_noise_pio_s1_chipselect),                               //                                                       .chipselect
		.onchip_memory2_0_s1_address                                  (mm_interconnect_0_onchip_memory2_0_s1_address),                           //                                    onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                    (mm_interconnect_0_onchip_memory2_0_s1_write),                             //                                                       .write
		.onchip_memory2_0_s1_readdata                                 (mm_interconnect_0_onchip_memory2_0_s1_readdata),                          //                                                       .readdata
		.onchip_memory2_0_s1_writedata                                (mm_interconnect_0_onchip_memory2_0_s1_writedata),                         //                                                       .writedata
		.onchip_memory2_0_s1_byteenable                               (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                        //                                                       .byteenable
		.onchip_memory2_0_s1_chipselect                               (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                        //                                                       .chipselect
		.onchip_memory2_0_s1_clken                                    (mm_interconnect_0_onchip_memory2_0_s1_clken),                             //                                                       .clken
		.piece_pio_s1_address                                         (mm_interconnect_0_piece_pio_s1_address),                                  //                                           piece_pio_s1.address
		.piece_pio_s1_write                                           (mm_interconnect_0_piece_pio_s1_write),                                    //                                                       .write
		.piece_pio_s1_readdata                                        (mm_interconnect_0_piece_pio_s1_readdata),                                 //                                                       .readdata
		.piece_pio_s1_writedata                                       (mm_interconnect_0_piece_pio_s1_writedata),                                //                                                       .writedata
		.piece_pio_s1_chipselect                                      (mm_interconnect_0_piece_pio_s1_chipselect),                               //                                                       .chipselect
		.sdram_s1_address                                             (mm_interconnect_0_sdram_s1_address),                                      //                                               sdram_s1.address
		.sdram_s1_write                                               (mm_interconnect_0_sdram_s1_write),                                        //                                                       .write
		.sdram_s1_read                                                (mm_interconnect_0_sdram_s1_read),                                         //                                                       .read
		.sdram_s1_readdata                                            (mm_interconnect_0_sdram_s1_readdata),                                     //                                                       .readdata
		.sdram_s1_writedata                                           (mm_interconnect_0_sdram_s1_writedata),                                    //                                                       .writedata
		.sdram_s1_byteenable                                          (mm_interconnect_0_sdram_s1_byteenable),                                   //                                                       .byteenable
		.sdram_s1_readdatavalid                                       (mm_interconnect_0_sdram_s1_readdatavalid),                                //                                                       .readdatavalid
		.sdram_s1_waitrequest                                         (mm_interconnect_0_sdram_s1_waitrequest),                                  //                                                       .waitrequest
		.sdram_s1_chipselect                                          (mm_interconnect_0_sdram_s1_chipselect),                                   //                                                       .chipselect
		.spi_0_spi_control_port_address                               (mm_interconnect_0_spi_0_spi_control_port_address),                        //                                 spi_0_spi_control_port.address
		.spi_0_spi_control_port_write                                 (mm_interconnect_0_spi_0_spi_control_port_write),                          //                                                       .write
		.spi_0_spi_control_port_read                                  (mm_interconnect_0_spi_0_spi_control_port_read),                           //                                                       .read
		.spi_0_spi_control_port_readdata                              (mm_interconnect_0_spi_0_spi_control_port_readdata),                       //                                                       .readdata
		.spi_0_spi_control_port_writedata                             (mm_interconnect_0_spi_0_spi_control_port_writedata),                      //                                                       .writedata
		.spi_0_spi_control_port_chipselect                            (mm_interconnect_0_spi_0_spi_control_port_chipselect),                     //                                                       .chipselect
		.sysid_qsys_0_control_slave_address                           (mm_interconnect_0_sysid_qsys_0_control_slave_address),                    //                             sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                          (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),                   //                                                       .readdata
		.timer_s1_address                                             (mm_interconnect_0_timer_s1_address),                                      //                                               timer_s1.address
		.timer_s1_write                                               (mm_interconnect_0_timer_s1_write),                                        //                                                       .write
		.timer_s1_readdata                                            (mm_interconnect_0_timer_s1_readdata),                                     //                                                       .readdata
		.timer_s1_writedata                                           (mm_interconnect_0_timer_s1_writedata),                                    //                                                       .writedata
		.timer_s1_chipselect                                          (mm_interconnect_0_timer_s1_chipselect),                                   //                                                       .chipselect
		.usb_gpx_s1_address                                           (mm_interconnect_0_usb_gpx_s1_address),                                    //                                             usb_gpx_s1.address
		.usb_gpx_s1_readdata                                          (mm_interconnect_0_usb_gpx_s1_readdata),                                   //                                                       .readdata
		.usb_irq_s1_address                                           (mm_interconnect_0_usb_irq_s1_address),                                    //                                             usb_irq_s1.address
		.usb_irq_s1_readdata                                          (mm_interconnect_0_usb_irq_s1_readdata),                                   //                                                       .readdata
		.usb_rst_s1_address                                           (mm_interconnect_0_usb_rst_s1_address),                                    //                                             usb_rst_s1.address
		.usb_rst_s1_write                                             (mm_interconnect_0_usb_rst_s1_write),                                      //                                                       .write
		.usb_rst_s1_readdata                                          (mm_interconnect_0_usb_rst_s1_readdata),                                   //                                                       .readdata
		.usb_rst_s1_writedata                                         (mm_interconnect_0_usb_rst_s1_writedata),                                  //                                                       .writedata
		.usb_rst_s1_chipselect                                        (mm_interconnect_0_usb_rst_s1_chipselect),                                 //                                                       .chipselect
		.VGA_text_mode_controller_0_avalon_mm_slave_address           (mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_address),    //             VGA_text_mode_controller_0_avalon_mm_slave.address
		.VGA_text_mode_controller_0_avalon_mm_slave_write             (mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_write),      //                                                       .write
		.VGA_text_mode_controller_0_avalon_mm_slave_read              (mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_read),       //                                                       .read
		.VGA_text_mode_controller_0_avalon_mm_slave_readdata          (mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_readdata),   //                                                       .readdata
		.VGA_text_mode_controller_0_avalon_mm_slave_writedata         (mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_writedata),  //                                                       .writedata
		.VGA_text_mode_controller_0_avalon_mm_slave_byteenable        (mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_byteenable), //                                                       .byteenable
		.VGA_text_mode_controller_0_avalon_mm_slave_chipselect        (mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_chipselect)  //                                                       .chipselect
	);

	labfinalsoc_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
